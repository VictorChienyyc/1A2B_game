magic
tech scmos
timestamp 1712175754
<< metal1 >>
rect -730 2212 -622 2230
rect -441 2204 -333 2222
rect -106 2218 2 2236
rect 175 2210 283 2228
rect 783 2213 891 2231
rect 1081 2213 1189 2231
rect -493 1482 -480 1492
rect -493 1466 -481 1482
rect -568 1456 -481 1466
rect 1009 1471 1018 1492
rect 933 1456 1021 1471
rect -568 1454 -488 1456
rect -110 1437 -43 1447
rect -110 1420 -70 1437
rect -560 1382 -534 1383
rect -560 -220 -534 1364
rect -97 1304 -74 1420
rect -316 1297 -74 1304
rect -325 1289 -74 1297
rect -325 1286 -83 1289
rect -325 1264 -314 1286
rect -326 1256 -311 1264
rect -328 62 -311 1256
rect -33 205 86 218
rect 103 205 110 218
rect -46 204 110 205
rect 1132 142 1151 1371
rect 118 138 129 139
rect 181 138 193 139
rect 118 118 193 138
rect -325 0 -314 62
rect 118 58 129 118
rect 181 82 193 118
rect -328 -2 -311 0
rect -328 -5 -9 -2
rect -328 -6 -42 -5
rect -13 -6 -9 -5
rect 9 -6 15 -2
rect -229 -12 -28 -11
rect -229 -17 -1 -12
rect 471 -16 629 -13
rect 1128 -16 1154 142
rect -229 -18 -28 -17
rect -229 -27 -176 -18
rect 205 -21 1154 -16
rect 3 -26 10 -22
rect 43 -23 47 -22
rect 36 -26 47 -23
rect 59 -26 1154 -21
rect -552 -355 -534 -220
rect -202 -307 -176 -27
rect 36 -34 40 -26
rect 205 -28 1154 -26
rect 205 -39 1151 -28
rect 205 -47 1090 -39
rect 1132 -47 1151 -39
rect 471 -48 633 -47
rect 471 -54 629 -48
rect 30 -187 42 -126
rect 180 -187 192 -61
rect 29 -196 192 -187
rect 29 -197 191 -196
rect 30 -231 44 -197
rect -202 -355 -172 -307
rect -552 -367 -172 -355
rect -552 -369 -490 -367
rect 37 -1380 44 -231
rect 37 -1389 121 -1380
rect 37 -1390 44 -1389
rect 111 -1490 118 -1389
<< m2contact >>
rect -581 1454 -568 1466
rect 920 1456 933 1475
rect -43 1437 -31 1449
rect -560 1364 -534 1382
rect 1132 1371 1151 1381
rect -46 205 -33 218
rect 86 205 103 219
rect 181 47 194 82
rect 5 -6 9 -2
rect 10 -26 14 -22
rect 36 -38 40 -34
rect 180 -61 193 -51
<< metal2 >>
rect -1478 1475 -1471 1482
rect -1405 1475 -1400 1490
rect -1478 1470 -1400 1475
rect -1176 1468 -1170 1486
rect -1107 1468 -1102 1490
rect -1176 1462 -1098 1468
rect -876 1461 -870 1486
rect -808 1461 -802 1492
rect -877 1450 -802 1461
rect -643 1306 -628 1484
rect -577 1474 -572 1483
rect -581 1466 -568 1474
rect -560 1418 -533 1483
rect -276 1469 -269 1486
rect -205 1469 -201 1490
rect -276 1462 -201 1469
rect -276 1460 -269 1462
rect -43 1449 -34 1485
rect 22 1451 30 1485
rect 94 1451 98 1495
rect 21 1441 99 1451
rect 257 1444 268 1488
rect 622 1468 628 1484
rect 694 1468 701 1492
rect 622 1458 701 1468
rect 22 1440 30 1441
rect -560 1382 -534 1418
rect 37 1413 62 1441
rect 94 1440 98 1441
rect -45 1408 62 1413
rect -560 1363 -534 1364
rect -46 1399 62 1408
rect -46 1397 56 1399
rect -1491 1295 -1450 1299
rect -1456 1228 -1450 1295
rect -755 1283 -628 1306
rect -755 1280 -630 1283
rect -1486 1224 -1447 1228
rect -1493 997 -1454 999
rect -1493 995 -1451 997
rect -1457 927 -1451 995
rect -1486 923 -1447 927
rect -1491 695 -1452 699
rect -1459 630 -1453 695
rect -1484 626 -1445 630
rect -1459 625 -1453 626
rect -1491 395 -1448 399
rect -1454 329 -1448 395
rect -1485 325 -1446 329
rect -1486 -29 -1447 -25
rect -1459 -95 -1453 -29
rect -1492 -99 -1453 -95
rect -755 -448 -722 1280
rect -46 218 -34 1397
rect 257 1394 275 1444
rect 858 1420 866 1485
rect 922 1475 929 1486
rect 1157 1484 1166 1489
rect 979 1482 1003 1483
rect 944 1474 1003 1482
rect 979 1473 1003 1474
rect 260 1324 275 1394
rect 849 1335 873 1420
rect 994 1417 1000 1473
rect 1222 1465 1229 1487
rect 1293 1465 1300 1490
rect 1222 1455 1300 1465
rect 1222 1454 1229 1455
rect 1293 1452 1300 1455
rect 992 1397 1002 1417
rect 1132 1397 1166 1399
rect 992 1385 1166 1397
rect 995 1384 1166 1385
rect 1132 1381 1166 1384
rect 1151 1376 1166 1381
rect -7 1312 284 1324
rect 544 1320 874 1335
rect -7 1303 163 1312
rect 257 1311 268 1312
rect -46 12 -34 205
rect -4 124 16 1303
rect -66 6 -34 12
rect 5 -2 9 124
rect 87 9 103 205
rect 180 47 181 82
rect 544 78 554 1320
rect 1467 1297 1493 1299
rect 1459 1295 1493 1297
rect 1459 1228 1470 1295
rect 1459 1224 1496 1228
rect 1464 997 1490 998
rect 1455 994 1490 997
rect 1455 927 1466 994
rect 1455 924 1484 927
rect 1458 923 1484 924
rect 1464 696 1490 699
rect 1457 695 1490 696
rect 1457 627 1468 695
rect 1457 623 1489 627
rect 1465 398 1491 399
rect 1459 395 1491 398
rect 1459 329 1470 395
rect 1459 325 1488 329
rect 1466 97 1492 98
rect 1455 94 1492 97
rect 87 3 130 9
rect 87 2 103 3
rect 10 -150 14 -26
rect 69 -34 73 -33
rect 40 -38 73 -34
rect 69 -150 73 -38
rect 180 -51 192 47
rect 541 -25 556 78
rect 1455 28 1466 94
rect 1455 24 1490 28
rect 180 -63 192 -61
rect 544 -146 554 -25
rect -74 -162 19 -150
rect 53 -151 343 -150
rect 544 -151 549 -146
rect -74 -448 -62 -162
rect 53 -165 591 -151
rect -755 -467 -62 -448
rect -1493 -505 -1454 -501
rect 1465 -503 1491 -500
rect -1460 -572 -1454 -505
rect 1462 -504 1491 -503
rect -1484 -576 -1445 -572
rect 1462 -573 1473 -504
rect 1461 -577 1487 -573
rect -1491 -804 -1452 -800
rect -1461 -874 -1455 -804
rect 1459 -806 1491 -802
rect 1459 -871 1470 -806
rect -1487 -878 -1448 -874
rect 1459 -875 1486 -871
rect -1492 -1105 -1452 -1101
rect 1464 -1103 1490 -1100
rect -1458 -1171 -1452 -1105
rect 1460 -1104 1490 -1103
rect -1484 -1175 -1445 -1171
rect 1460 -1174 1471 -1104
rect 1460 -1176 1487 -1174
rect 1461 -1178 1487 -1176
rect -1482 -1401 -1475 -1400
rect -1491 -1405 -1475 -1401
rect 1469 -1402 1495 -1401
rect -1478 -1470 -1475 -1405
rect 1464 -1405 1495 -1402
rect -1105 -1420 -1099 -1419
rect -1178 -1430 -1099 -1420
rect -1482 -1471 -1401 -1470
rect -1482 -1476 -1399 -1471
rect -1482 -1483 -1468 -1476
rect -1405 -1490 -1399 -1476
rect -1178 -1484 -1170 -1430
rect -1105 -1491 -1099 -1430
rect -876 -1432 -870 -1423
rect -804 -1432 -798 -1428
rect -876 -1437 -798 -1432
rect -876 -1484 -870 -1437
rect -804 -1489 -798 -1437
rect -577 -1438 -499 -1429
rect 23 -1437 101 -1436
rect -577 -1485 -571 -1438
rect -505 -1490 -499 -1438
rect 22 -1443 101 -1437
rect 324 -1443 331 -1442
rect 22 -1485 31 -1443
rect 96 -1492 100 -1443
rect 324 -1449 403 -1443
rect 324 -1486 331 -1449
rect 396 -1490 403 -1449
rect 623 -1445 630 -1434
rect 696 -1445 703 -1440
rect 623 -1452 703 -1445
rect 623 -1485 630 -1452
rect 696 -1491 703 -1452
rect 923 -1451 929 -1447
rect 996 -1451 1002 -1450
rect 1224 -1451 1232 -1450
rect 923 -1461 1004 -1451
rect 1224 -1459 1303 -1451
rect 923 -1488 929 -1461
rect 996 -1491 1002 -1461
rect 1224 -1483 1232 -1459
rect 1295 -1492 1301 -1459
rect 1464 -1472 1475 -1405
rect 1462 -1476 1488 -1472
use PadFC  16_0
timestamp 1000338511
transform 1 0 -2500 0 1 1500
box 327 -3 1003 673
use PadFC  16_1
timestamp 1000338511
transform 0 1 1500 -1 0 2500
box 327 -3 1003 673
use PadFC  16_2
timestamp 1000338511
transform 0 -1 -1500 1 0 -2500
box 327 -3 1003 673
use PadFC  16_3
timestamp 1000338511
transform -1 0 2500 0 -1 -1500
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 1200
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 900
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 600
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 300
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 0
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -600
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -900
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1200
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 1500 1 0 1200
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 1500 1 0 900
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 1500 1 0 600
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 1500 1 0 300
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 1500 1 0 0
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 1500 1 0 -600
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 1500 1 0 -900
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 1500 1 0 -1200
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1500
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 1500 1 0 -1500
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1500
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 1500
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1500
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 300
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 1500 -1 0 0
box -3 -11 303 1000
use hwtest  hwtest_0
timestamp 1712112060
transform 1 0 -111 0 1 -149
box 14 13 266 227
<< labels >>
rlabel metal1 202 2220 202 2220 1 p_d
rlabel metal1 -85 2226 -85 2226 1 p_b
rlabel metal1 -419 2216 -419 2217 1 p_i
rlabel metal1 809 2223 809 2223 1 p_c
rlabel metal1 1124 2228 1124 2228 1 p_h
rlabel metal1 -704 2223 -704 2223 1 p_a
rlabel metal1 -19 -3 -19 -3 1 b
rlabel metal1 -14 -15 -14 -15 1 i
rlabel metal2 12 -89 12 -89 1 a
rlabel metal2 7 1 7 1 1 d
rlabel metal2 71 -89 71 -89 1 c
rlabel metal1 61 -24 61 -24 1 h
rlabel metal1 203 -23 203 -23 1 h
rlabel metal1 233 -35 233 -35 1 j
<< end >>
