magic
tech scmos
magscale 1 2
timestamp 1714524297
<< metal1 >>
rect 28 3614 3796 3654
rect 76 3566 3748 3606
rect 76 3534 3748 3546
rect 757 3467 1144 3473
rect 1797 3467 1848 3473
rect 1973 3467 2120 3473
rect 2741 3467 2792 3473
rect 2901 3467 3048 3473
rect 1045 3447 1160 3453
rect 1221 3447 1240 3453
rect 1749 3447 1784 3453
rect 2197 3447 2216 3453
rect 2728 3447 2808 3453
rect 2869 3447 2888 3453
rect 3064 3447 3096 3453
rect 3157 3447 3240 3453
rect 1592 3427 1611 3433
rect 28 3334 3796 3346
rect 1477 3267 1512 3273
rect 1480 3247 1499 3253
rect 693 3227 776 3233
rect 1013 3227 1032 3233
rect 1240 3227 1259 3233
rect 1432 3232 1467 3233
rect 1432 3227 1496 3232
rect 1637 3227 1720 3233
rect 2104 3227 2155 3233
rect 2216 3227 2235 3233
rect 2248 3227 2267 3233
rect 2328 3227 2379 3233
rect 2488 3227 2523 3233
rect 2600 3227 2619 3233
rect 2632 3227 2651 3233
rect 3048 3227 3099 3233
rect 693 3207 760 3213
rect 824 3207 859 3213
rect 1253 3210 1259 3227
rect 1461 3226 1496 3227
rect 1333 3207 1368 3213
rect 1832 3207 1851 3213
rect 2229 3210 2235 3227
rect 2261 3210 2267 3227
rect 2373 3190 2379 3227
rect 2613 3210 2619 3227
rect 2645 3210 2651 3227
rect 76 3134 3748 3146
rect 421 3051 427 3073
rect 1029 3053 1035 3070
rect 1573 3053 1579 3070
rect 1845 3053 1851 3070
rect 2485 3053 2491 3090
rect 2517 3067 2536 3073
rect 565 3047 600 3053
rect 725 3047 744 3053
rect 1016 3047 1035 3053
rect 1077 3013 1083 3050
rect 1416 3047 1467 3053
rect 1528 3047 1579 3053
rect 1688 3047 1739 3053
rect 1800 3047 1851 3053
rect 1864 3047 1899 3053
rect 1941 3047 1992 3053
rect 2168 3047 2219 3053
rect 2440 3047 2491 3053
rect 2520 3047 2539 3053
rect 2645 3047 2680 3053
rect 3032 3047 3083 3053
rect 3157 3047 3192 3053
rect 3253 3047 3304 3053
rect 421 3007 440 3013
rect 1061 3007 1083 3013
rect 28 2934 3796 2946
rect 421 2833 427 2853
rect 421 2827 555 2833
rect 773 2813 779 2853
rect 1864 2847 1883 2853
rect 1144 2827 1195 2833
rect 1320 2827 1371 2833
rect 1432 2827 1483 2833
rect 1496 2827 1531 2833
rect 1592 2827 1643 2833
rect 1656 2827 1752 2833
rect 1813 2827 1832 2833
rect 1861 2827 1896 2833
rect 2104 2827 2155 2833
rect 2600 2827 2651 2833
rect 2712 2827 2763 2833
rect 2872 2827 2923 2833
rect 3016 2827 3048 2833
rect 3109 2827 3128 2833
rect 3221 2827 3272 2833
rect 3333 2827 3368 2833
rect 773 2807 856 2813
rect 1208 2807 1227 2813
rect 1352 2807 1368 2813
rect 1509 2807 1528 2813
rect 1637 2810 1643 2827
rect 1784 2807 1803 2813
rect 2296 2807 2312 2813
rect 2757 2790 2763 2827
rect 3157 2807 3256 2813
rect 76 2734 3748 2746
rect 869 2654 875 2670
rect 1208 2667 1227 2673
rect 552 2647 587 2653
rect 856 2648 875 2654
rect 997 2653 1032 2654
rect 1349 2653 1355 2690
rect 1720 2667 1739 2673
rect 1784 2667 1819 2673
rect 1893 2667 1960 2673
rect 2213 2653 2219 2690
rect 2245 2667 2264 2673
rect 2757 2653 2763 2690
rect 2789 2667 2808 2673
rect 3109 2654 3115 2670
rect 3333 2654 3339 2670
rect 968 2648 1032 2653
rect 968 2647 1003 2648
rect 1144 2647 1195 2653
rect 1304 2647 1355 2653
rect 1688 2647 1723 2653
rect 1813 2647 1832 2653
rect 1896 2647 1931 2653
rect 1976 2647 1995 2653
rect 2168 2647 2219 2653
rect 2248 2647 2267 2653
rect 2520 2647 2539 2653
rect 2712 2647 2763 2653
rect 2792 2647 2811 2653
rect 2984 2647 3035 2653
rect 3096 2648 3115 2654
rect 3208 2647 3259 2653
rect 3320 2648 3339 2654
rect 28 2534 3796 2546
rect 600 2427 683 2433
rect 981 2427 1032 2433
rect 1272 2427 1339 2433
rect 1400 2427 1451 2433
rect 1624 2427 1675 2433
rect 1829 2413 1835 2429
rect 1925 2427 1976 2433
rect 2184 2427 2235 2433
rect 2264 2427 2283 2433
rect 2472 2427 2523 2433
rect 2552 2427 2571 2433
rect 2760 2427 2779 2433
rect 613 2407 680 2413
rect 981 2407 1016 2413
rect 1157 2407 1208 2413
rect 1317 2407 1336 2413
rect 1464 2407 1483 2413
rect 1688 2407 1835 2413
rect 1880 2407 1963 2413
rect 2024 2407 2107 2413
rect 1477 2393 1483 2407
rect 1477 2387 1547 2393
rect 2229 2390 2235 2427
rect 2261 2407 2280 2413
rect 2389 2407 2408 2413
rect 2389 2387 2395 2407
rect 2517 2390 2523 2427
rect 2901 2413 2907 2433
rect 2965 2427 3016 2433
rect 3077 2427 3096 2433
rect 2549 2407 2568 2413
rect 2664 2407 2699 2413
rect 2725 2407 2744 2413
rect 2757 2407 2776 2413
rect 2872 2407 2907 2413
rect 2949 2407 3000 2413
rect 2693 2387 2728 2393
rect 76 2334 3748 2346
rect 789 2253 795 2270
rect 821 2267 888 2273
rect 1253 2267 1304 2273
rect 1560 2267 1627 2273
rect 981 2253 1016 2254
rect 1861 2253 1867 2290
rect 1880 2267 1899 2273
rect 2165 2267 2344 2273
rect 2629 2267 2712 2273
rect 3016 2267 3035 2273
rect 3253 2254 3259 2270
rect 776 2247 795 2253
rect 952 2248 1016 2253
rect 952 2247 987 2248
rect 1205 2247 1240 2253
rect 1368 2247 1419 2253
rect 1496 2247 1547 2253
rect 1704 2247 1755 2253
rect 1816 2247 1867 2253
rect 2008 2247 2027 2253
rect 2133 2247 2152 2253
rect 2936 2247 2955 2253
rect 3240 2248 3259 2254
rect 1000 2227 1019 2233
rect 28 2134 3796 2146
rect 664 2027 683 2033
rect 856 2027 875 2033
rect 1208 2027 1259 2033
rect 1333 2027 1352 2033
rect 1432 2027 1483 2033
rect 1637 2027 1656 2033
rect 1736 2027 1787 2033
rect 1848 2027 1899 2033
rect 2328 2027 2347 2033
rect 2456 2027 2507 2033
rect 2536 2027 2555 2033
rect 2728 2027 2779 2033
rect 1893 1990 1899 2027
rect 1912 2007 1963 2013
rect 1973 2007 1992 2013
rect 2341 2010 2347 2027
rect 2373 2007 2392 2013
rect 1973 1993 1979 2007
rect 1925 1987 1979 1993
rect 2501 1990 2507 2027
rect 2840 2026 2859 2032
rect 2872 2027 2952 2033
rect 3013 2027 3064 2033
rect 3077 2027 3224 2033
rect 2533 2007 2552 2013
rect 2853 2010 2859 2026
rect 2917 2007 2936 2013
rect 3237 2007 3272 2013
rect 76 1934 3748 1946
rect 1237 1867 1288 1873
rect 1352 1867 1435 1873
rect 1685 1853 1691 1869
rect 1717 1854 1723 1869
rect 2165 1867 2232 1873
rect 616 1847 651 1853
rect 917 1847 952 1853
rect 965 1847 984 1853
rect 1112 1847 1147 1853
rect 1285 1847 1304 1853
rect 1512 1847 1563 1853
rect 1624 1847 1691 1853
rect 1704 1848 1723 1854
rect 2261 1853 2267 1869
rect 1797 1847 1944 1853
rect 2024 1847 2059 1853
rect 2248 1847 2267 1853
rect 2312 1847 2347 1853
rect 2389 1847 2440 1853
rect 2501 1847 2507 1869
rect 2885 1854 2891 1869
rect 2872 1848 2891 1854
rect 3221 1853 3227 1869
rect 3253 1867 3272 1873
rect 3480 1867 3499 1873
rect 2904 1847 2923 1853
rect 3064 1847 3115 1853
rect 3176 1847 3227 1853
rect 3240 1847 3259 1853
rect 3397 1847 3416 1853
rect 28 1734 3796 1746
rect 1016 1647 1115 1653
rect 584 1627 603 1633
rect 616 1627 664 1633
rect 693 1627 840 1633
rect 888 1627 984 1633
rect 1176 1626 1195 1632
rect 1352 1627 1403 1633
rect 1557 1627 1576 1633
rect 1704 1626 1723 1632
rect 1989 1627 2008 1633
rect 2101 1627 2120 1633
rect 2181 1627 2232 1633
rect 2293 1627 2312 1633
rect 2357 1627 2456 1633
rect 2469 1627 2488 1633
rect 2744 1627 2763 1633
rect 2904 1627 2955 1633
rect 696 1607 731 1613
rect 853 1607 872 1613
rect 1016 1607 1131 1613
rect 1189 1610 1195 1626
rect 1256 1607 1275 1613
rect 1717 1610 1723 1626
rect 2389 1607 2440 1613
rect 2757 1610 2763 1627
rect 3269 1613 3275 1629
rect 3397 1627 3416 1633
rect 3205 1607 3256 1613
rect 3269 1607 3304 1613
rect 3157 1587 3240 1593
rect 76 1534 3748 1546
rect 485 1487 600 1493
rect 597 1467 760 1473
rect 789 1467 808 1473
rect 933 1467 952 1473
rect 981 1467 1016 1473
rect 1045 1467 1064 1473
rect 1112 1467 1195 1473
rect 1589 1467 1608 1473
rect 1589 1453 1595 1467
rect 2549 1453 2555 1490
rect 2581 1467 2600 1473
rect 3336 1467 3355 1473
rect 3397 1467 3496 1473
rect 805 1447 824 1453
rect 968 1447 1019 1453
rect 1032 1447 1080 1453
rect 1413 1447 1448 1453
rect 1573 1447 1595 1453
rect 1672 1447 1723 1453
rect 1925 1447 1992 1453
rect 2504 1447 2555 1453
rect 2584 1447 2603 1453
rect 3112 1447 3163 1453
rect 3237 1447 3272 1453
rect 3336 1447 3384 1453
rect 1717 1433 1723 1447
rect 1717 1427 1752 1433
rect 28 1334 3796 1346
rect 917 1267 955 1273
rect 885 1247 936 1253
rect 485 1227 536 1233
rect 648 1227 667 1233
rect 728 1227 827 1233
rect 949 1230 955 1267
rect 984 1247 1003 1253
rect 1576 1247 1659 1253
rect 2136 1247 2155 1253
rect 3416 1247 3435 1253
rect 1560 1227 1595 1233
rect 549 1207 600 1213
rect 661 1193 667 1227
rect 1688 1226 1707 1232
rect 677 1207 696 1213
rect 789 1207 824 1213
rect 1013 1207 1096 1213
rect 1109 1207 1240 1213
rect 1573 1207 1672 1213
rect 1701 1211 1707 1226
rect 1989 1211 1995 1233
rect 2120 1227 2219 1233
rect 2293 1227 2328 1233
rect 2408 1227 2427 1233
rect 2600 1227 2651 1233
rect 2725 1227 2744 1233
rect 3445 1227 3464 1233
rect 3544 1227 3579 1233
rect 2133 1207 2216 1213
rect 3096 1207 3128 1213
rect 3304 1207 3323 1213
rect 3557 1207 3576 1213
rect 661 1187 680 1193
rect 76 1134 3748 1146
rect 837 1087 904 1093
rect 805 1067 920 1073
rect 1045 1067 1064 1073
rect 1125 1067 1144 1073
rect 392 1047 443 1053
rect 517 1047 536 1053
rect 805 1047 811 1067
rect 1189 1047 1195 1069
rect 1221 1067 1256 1073
rect 1608 1067 1675 1073
rect 1957 1067 2008 1073
rect 1253 1047 1272 1053
rect 1301 1047 1336 1053
rect 1605 1047 1720 1053
rect 1781 1047 1800 1053
rect 1893 1047 1944 1053
rect 2037 1047 2043 1069
rect 2133 1053 2139 1069
rect 2213 1053 2219 1069
rect 3349 1067 3366 1073
rect 3397 1067 3480 1073
rect 3349 1053 3355 1067
rect 3509 1053 3515 1069
rect 2133 1047 2219 1053
rect 2408 1047 2427 1053
rect 2661 1047 2680 1053
rect 2824 1047 2859 1053
rect 3016 1047 3067 1053
rect 3338 1047 3355 1053
rect 3384 1047 3467 1053
rect 3496 1047 3515 1053
rect 3576 1047 3611 1053
rect 792 1027 827 1033
rect 1192 1027 1211 1033
rect 1413 1027 1448 1033
rect 28 934 3796 946
rect 997 867 1099 873
rect 613 847 635 853
rect 664 847 699 853
rect 997 847 1080 853
rect 613 833 619 847
rect 693 833 699 847
rect 552 827 619 833
rect 629 827 648 833
rect 693 827 712 833
rect 773 827 792 833
rect 984 827 1019 833
rect 1093 830 1099 867
rect 1128 847 1243 853
rect 1608 847 1659 853
rect 1141 827 1272 833
rect 1333 827 1416 833
rect 1461 827 1579 833
rect 1592 827 1643 833
rect 1944 827 1995 833
rect 2088 827 2155 833
rect 2232 827 2283 833
rect 2357 827 2376 833
rect 2504 827 2587 833
rect 2776 827 2827 833
rect 3032 827 3083 833
rect 3397 827 3496 833
rect 3560 827 3611 833
rect 517 807 536 813
rect 549 807 632 813
rect 757 807 776 813
rect 805 807 904 813
rect 1173 807 1256 813
rect 1285 807 1304 813
rect 1349 807 1400 813
rect 1448 807 1563 813
rect 1573 810 1579 827
rect 2421 807 2456 813
rect 2488 807 2507 813
rect 2581 810 2587 827
rect 2680 807 2699 813
rect 3336 807 3355 813
rect 3560 807 3579 813
rect 757 790 763 807
rect 2421 767 2427 807
rect 76 734 3748 746
rect 517 667 536 673
rect 549 667 568 673
rect 597 667 680 673
rect 725 653 731 670
rect 392 647 443 653
rect 504 647 523 653
rect 552 647 584 653
rect 629 647 696 653
rect 725 647 747 653
rect 901 651 907 673
rect 949 667 968 673
rect 1224 667 1243 673
rect 1813 667 1912 673
rect 2085 667 2104 673
rect 2501 667 2520 673
rect 2629 667 2648 673
rect 2744 667 2763 673
rect 2853 667 2888 673
rect 3208 667 3227 673
rect 3333 667 3352 673
rect 3448 667 3512 673
rect 3557 653 3563 670
rect 1221 647 1320 653
rect 1365 647 1400 653
rect 1496 647 1515 653
rect 1800 647 1883 653
rect 1960 647 1979 653
rect 1989 647 2072 653
rect 2165 647 2248 653
rect 2277 647 2328 653
rect 2405 647 2440 653
rect 2485 647 2536 653
rect 2616 647 2651 653
rect 2920 647 2939 653
rect 3320 647 3355 653
rect 3496 647 3515 653
rect 3557 647 3579 653
rect 1973 633 1979 647
rect 888 627 907 633
rect 1045 627 1112 633
rect 1973 627 2027 633
rect 789 607 920 613
rect 28 534 3796 546
rect 2712 447 2811 453
rect 3160 447 3243 453
rect 728 427 747 433
rect 1224 427 1243 433
rect 1493 413 1499 429
rect 1509 427 1528 433
rect 1589 427 1640 433
rect 1912 427 1963 433
rect 2037 427 2056 433
rect 2085 427 2200 433
rect 2344 427 2379 433
rect 2565 427 2648 433
rect 2661 427 2680 433
rect 2773 427 2824 433
rect 2888 427 2923 433
rect 3013 427 3096 433
rect 3109 427 3128 433
rect 3157 427 3256 433
rect 3333 427 3368 433
rect 3381 427 3432 433
rect 3496 427 3531 433
rect 1381 407 1464 413
rect 1493 407 1512 413
rect 1541 407 1624 413
rect 2357 407 2376 413
rect 2472 407 2507 413
rect 2520 407 2619 413
rect 2712 407 2747 413
rect 2901 407 2920 413
rect 3016 407 3051 413
rect 3509 407 3528 413
rect 2501 390 2507 407
rect 2613 387 2619 407
rect 76 334 3748 346
rect 1733 273 1739 290
rect 2981 287 3032 293
rect 1525 267 1576 273
rect 1589 267 1704 273
rect 1733 267 1752 273
rect 2293 253 2299 273
rect 2501 253 2507 273
rect 2949 253 2955 270
rect 1208 247 1259 253
rect 1333 247 1352 253
rect 1592 247 1688 253
rect 1749 247 1768 253
rect 2293 247 2552 253
rect 2696 247 2731 253
rect 2837 247 2856 253
rect 2920 247 2955 253
rect 3077 247 3240 253
rect 1464 227 1483 233
rect 28 134 3796 146
rect 76 74 3748 114
rect 28 26 3796 66
<< metal2 >>
rect 28 26 68 3654
rect 76 74 116 3606
rect 693 3253 699 3273
rect 357 3087 395 3093
rect 357 3067 363 3087
rect 405 3027 411 3253
rect 613 3227 619 3253
rect 661 3247 699 3253
rect 549 3187 555 3213
rect 645 3173 651 3213
rect 661 3207 667 3247
rect 677 3187 683 3233
rect 693 3227 699 3247
rect 709 3213 715 3233
rect 693 3207 715 3213
rect 693 3173 699 3207
rect 645 3167 699 3173
rect 421 3067 427 3113
rect 453 3027 459 3093
rect 469 3013 475 3073
rect 565 3067 571 3113
rect 565 3013 571 3053
rect 421 2847 427 3013
rect 469 3007 571 3013
rect 581 2873 587 3073
rect 613 2933 619 3053
rect 725 3027 731 3053
rect 757 2993 763 3473
rect 789 3107 795 3213
rect 805 3147 811 3233
rect 789 3067 811 3073
rect 741 2987 763 2993
rect 613 2927 651 2933
rect 549 2867 587 2873
rect 549 2827 555 2867
rect 517 2807 555 2813
rect 645 2807 651 2927
rect 741 2833 747 2987
rect 741 2827 763 2833
rect 773 2827 779 3053
rect 805 3027 811 3053
rect 821 2933 827 3493
rect 1125 3487 1179 3493
rect 965 3247 1019 3253
rect 917 3227 939 3233
rect 837 3113 843 3173
rect 853 3133 859 3213
rect 869 3173 875 3213
rect 965 3207 971 3247
rect 981 3187 987 3213
rect 997 3173 1003 3233
rect 1013 3227 1019 3247
rect 869 3167 1003 3173
rect 1013 3147 1019 3213
rect 1045 3173 1051 3453
rect 1125 3227 1131 3487
rect 1141 3447 1147 3473
rect 1173 3467 1179 3487
rect 1205 3467 1211 3493
rect 1477 3467 1483 3573
rect 1605 3453 1611 3493
rect 1189 3447 1227 3453
rect 1589 3447 1611 3453
rect 1477 3267 1483 3373
rect 1589 3333 1595 3447
rect 1605 3407 1611 3433
rect 1637 3427 1643 3573
rect 1653 3413 1659 3473
rect 1749 3467 1755 3493
rect 1765 3467 1803 3473
rect 1749 3413 1755 3453
rect 1621 3373 1627 3413
rect 1653 3407 1755 3413
rect 1765 3373 1771 3467
rect 1621 3367 1771 3373
rect 1589 3327 1643 3333
rect 1493 3287 1611 3293
rect 1493 3247 1499 3287
rect 1525 3247 1531 3273
rect 1077 3187 1083 3213
rect 1045 3167 1083 3173
rect 853 3127 939 3133
rect 837 3107 859 3113
rect 805 2927 827 2933
rect 549 2747 555 2807
rect 757 2787 763 2827
rect 805 2793 811 2927
rect 853 2913 859 3107
rect 901 3047 907 3073
rect 933 3033 939 3127
rect 1029 3067 1035 3093
rect 789 2787 811 2793
rect 837 2907 859 2913
rect 917 3027 939 3033
rect 997 3047 1051 3053
rect 581 2647 587 2673
rect 597 2473 603 2773
rect 789 2753 795 2787
rect 837 2753 843 2907
rect 917 2893 923 3027
rect 997 2973 1003 3047
rect 1061 3027 1067 3053
rect 1061 2987 1067 3013
rect 773 2747 795 2753
rect 829 2747 843 2753
rect 853 2887 923 2893
rect 965 2967 1003 2973
rect 629 2727 747 2733
rect 629 2667 635 2727
rect 613 2627 619 2653
rect 645 2647 651 2673
rect 661 2573 667 2673
rect 693 2587 699 2673
rect 741 2647 747 2727
rect 773 2573 779 2747
rect 829 2613 835 2747
rect 821 2607 835 2613
rect 821 2573 827 2607
rect 853 2593 859 2887
rect 917 2827 923 2873
rect 949 2767 955 2813
rect 965 2807 971 2967
rect 1029 2827 1035 2853
rect 1061 2773 1067 2813
rect 869 2667 875 2693
rect 885 2627 891 2653
rect 853 2587 875 2593
rect 661 2567 779 2573
rect 805 2567 827 2573
rect 597 2467 619 2473
rect 613 2333 619 2467
rect 677 2447 731 2453
rect 677 2427 683 2447
rect 693 2427 715 2433
rect 725 2427 731 2447
rect 709 2407 731 2413
rect 565 2327 619 2333
rect 741 2333 747 2567
rect 741 2327 763 2333
rect 565 2213 571 2327
rect 613 2267 619 2313
rect 565 2207 587 2213
rect 581 2007 587 2207
rect 661 1993 667 2253
rect 757 2173 763 2327
rect 805 2293 811 2567
rect 853 2407 859 2433
rect 869 2387 875 2587
rect 901 2513 907 2713
rect 997 2667 1003 2693
rect 1013 2653 1019 2773
rect 1045 2767 1067 2773
rect 1045 2707 1051 2767
rect 893 2507 907 2513
rect 997 2647 1019 2653
rect 893 2373 899 2507
rect 965 2413 971 2433
rect 981 2427 987 2453
rect 965 2407 987 2413
rect 893 2367 907 2373
rect 901 2327 907 2367
rect 965 2347 971 2407
rect 997 2373 1003 2647
rect 1013 2607 1019 2633
rect 1029 2453 1035 2693
rect 1061 2627 1067 2753
rect 1077 2667 1083 3167
rect 1109 3027 1115 3153
rect 1125 3067 1131 3093
rect 1093 2927 1099 3013
rect 1189 2987 1195 3053
rect 1221 2987 1227 3073
rect 1237 3067 1243 3233
rect 1253 3227 1275 3233
rect 1605 3227 1611 3287
rect 1637 3227 1643 3327
rect 1333 3087 1339 3213
rect 1461 3173 1467 3213
rect 1445 3167 1467 3173
rect 1285 3047 1307 3053
rect 1333 3027 1339 3073
rect 1349 3067 1355 3113
rect 1173 2687 1179 2833
rect 1189 2827 1227 2833
rect 1189 2787 1195 2813
rect 1221 2787 1227 2813
rect 1237 2773 1243 2873
rect 1189 2767 1243 2773
rect 1189 2687 1195 2767
rect 1045 2607 1067 2613
rect 1093 2607 1115 2613
rect 1061 2487 1067 2607
rect 1029 2447 1051 2453
rect 1045 2413 1051 2447
rect 1109 2427 1115 2607
rect 1173 2533 1179 2673
rect 1221 2667 1227 2733
rect 1253 2707 1259 2813
rect 1349 2807 1355 3053
rect 1445 2887 1451 3167
rect 1541 3153 1547 3213
rect 1461 3067 1467 3153
rect 1541 3147 1611 3153
rect 1461 3007 1467 3053
rect 1365 2827 1371 2873
rect 1477 2847 1515 2853
rect 1477 2827 1483 2847
rect 1365 2793 1371 2813
rect 1349 2787 1371 2793
rect 1189 2647 1227 2653
rect 1237 2627 1243 2693
rect 1333 2667 1339 2773
rect 1205 2533 1211 2613
rect 1349 2587 1355 2787
rect 1461 2767 1467 2813
rect 1477 2733 1483 2813
rect 1509 2807 1515 2833
rect 1525 2827 1531 2853
rect 1557 2827 1563 3133
rect 1605 3113 1611 3147
rect 1637 3127 1643 3213
rect 1701 3187 1707 3213
rect 1717 3113 1723 3333
rect 1765 3293 1771 3367
rect 1765 3287 1787 3293
rect 1781 3227 1787 3287
rect 1797 3273 1803 3433
rect 1941 3407 1947 3473
rect 1973 3447 1979 3473
rect 2133 3413 2139 3453
rect 2117 3407 2139 3413
rect 2117 3313 2123 3407
rect 1797 3267 1835 3273
rect 1733 3147 1739 3213
rect 1829 3153 1835 3267
rect 1845 3227 1851 3253
rect 1845 3173 1851 3213
rect 1861 3207 1867 3313
rect 2005 3307 2027 3313
rect 2117 3307 2139 3313
rect 1893 3267 1979 3273
rect 1877 3187 1883 3233
rect 1893 3173 1899 3267
rect 1909 3247 1931 3253
rect 1845 3167 1899 3173
rect 1829 3147 1851 3153
rect 1605 3107 1739 3113
rect 1589 3047 1595 3073
rect 1605 3053 1611 3107
rect 1621 3067 1627 3093
rect 1605 3047 1627 3053
rect 1605 3007 1611 3033
rect 1381 2727 1483 2733
rect 1365 2627 1371 2673
rect 1381 2667 1387 2727
rect 1397 2667 1403 2713
rect 1493 2687 1514 2693
rect 1173 2527 1211 2533
rect 981 2367 1003 2373
rect 1029 2407 1051 2413
rect 805 2287 843 2293
rect 789 2267 827 2273
rect 741 2167 763 2173
rect 805 2247 827 2253
rect 677 2047 731 2053
rect 677 2027 683 2047
rect 693 2027 715 2033
rect 725 2027 731 2047
rect 677 2007 699 2013
rect 709 1993 715 2013
rect 741 2007 747 2167
rect 805 2027 811 2247
rect 837 2147 843 2287
rect 981 2167 987 2367
rect 1029 2307 1035 2407
rect 1013 2207 1019 2233
rect 1045 2227 1051 2393
rect 1141 2347 1147 2413
rect 1157 2407 1163 2453
rect 1109 2213 1115 2293
rect 1205 2267 1211 2527
rect 1381 2473 1387 2653
rect 1445 2647 1467 2653
rect 1493 2607 1499 2673
rect 1508 2667 1514 2687
rect 1333 2467 1387 2473
rect 1301 2313 1307 2413
rect 1317 2407 1323 2453
rect 1333 2427 1339 2467
rect 1285 2307 1307 2313
rect 1221 2267 1227 2293
rect 869 2047 923 2053
rect 869 2027 875 2047
rect 885 2027 907 2033
rect 917 2027 923 2047
rect 853 2007 875 2013
rect 661 1987 715 1993
rect 901 1967 907 2013
rect 933 1913 939 2053
rect 917 1907 939 1913
rect 597 1847 603 1873
rect 677 1867 683 1893
rect 629 1693 635 1833
rect 645 1813 651 1853
rect 725 1813 731 1853
rect 821 1847 843 1853
rect 917 1847 923 1907
rect 965 1893 971 2153
rect 1029 2067 1035 2213
rect 1109 2207 1131 2213
rect 1173 2207 1179 2253
rect 1013 1967 1019 2033
rect 1125 2027 1131 2207
rect 1205 2027 1211 2253
rect 1253 2247 1259 2293
rect 1221 2133 1227 2173
rect 1285 2133 1291 2307
rect 1221 2127 1235 2133
rect 1285 2127 1307 2133
rect 1229 2013 1235 2127
rect 1157 1907 1163 2013
rect 1221 2007 1235 2013
rect 965 1887 1035 1893
rect 933 1833 939 1873
rect 965 1867 1003 1873
rect 965 1833 971 1853
rect 933 1827 971 1833
rect 645 1807 667 1813
rect 725 1807 747 1813
rect 661 1773 667 1807
rect 661 1767 699 1773
rect 597 1687 635 1693
rect 565 1607 571 1633
rect 597 1627 603 1687
rect 629 1627 635 1653
rect 693 1647 699 1767
rect 741 1673 747 1807
rect 997 1793 1003 1867
rect 725 1667 747 1673
rect 981 1787 1003 1793
rect 645 1627 699 1633
rect 485 1193 491 1493
rect 597 1467 603 1613
rect 645 1607 651 1627
rect 725 1607 731 1667
rect 981 1653 987 1787
rect 1029 1673 1035 1887
rect 1061 1867 1067 1893
rect 1029 1667 1051 1673
rect 629 1373 635 1453
rect 741 1427 747 1453
rect 757 1393 763 1633
rect 821 1607 859 1613
rect 853 1587 859 1607
rect 901 1527 907 1653
rect 981 1647 1003 1653
rect 997 1613 1003 1647
rect 789 1487 827 1493
rect 773 1467 795 1473
rect 613 1367 635 1373
rect 741 1387 763 1393
rect 477 1187 491 1193
rect 517 1207 555 1213
rect 341 587 347 1073
rect 437 1047 443 1113
rect 477 1053 483 1187
rect 517 1153 523 1207
rect 501 1147 523 1153
rect 477 1047 491 1053
rect 485 1013 491 1047
rect 501 1027 507 1147
rect 517 1067 555 1073
rect 565 1067 571 1113
rect 549 1053 555 1067
rect 517 1013 523 1053
rect 549 1047 603 1053
rect 485 1007 523 1013
rect 453 847 459 933
rect 469 787 475 833
rect 485 813 491 873
rect 565 853 571 1033
rect 501 847 571 853
rect 485 807 523 813
rect 549 793 555 813
rect 517 787 555 793
rect 437 727 491 733
rect 437 647 443 727
rect 485 673 491 727
rect 597 693 603 1047
rect 613 1033 619 1367
rect 741 1233 747 1387
rect 741 1227 763 1233
rect 661 1207 683 1213
rect 661 1073 667 1207
rect 677 1093 683 1193
rect 677 1087 699 1093
rect 661 1067 683 1073
rect 613 1027 635 1033
rect 629 893 635 1027
rect 613 887 635 893
rect 613 833 619 887
rect 677 873 683 1067
rect 693 1047 699 1087
rect 725 1047 731 1073
rect 741 1067 747 1093
rect 757 1047 763 1227
rect 789 1207 795 1453
rect 805 1427 811 1453
rect 821 1227 827 1487
rect 869 1247 875 1353
rect 837 1087 843 1233
rect 869 1187 875 1213
rect 789 1033 795 1073
rect 725 993 731 1033
rect 717 987 731 993
rect 741 1027 795 1033
rect 677 867 699 873
rect 629 847 667 853
rect 613 827 635 833
rect 517 687 603 693
rect 485 667 523 673
rect 549 653 555 673
rect 597 667 603 687
rect 517 647 555 653
rect 629 647 635 813
rect 661 747 667 847
rect 693 733 699 867
rect 717 853 723 987
rect 717 847 731 853
rect 725 767 731 847
rect 741 813 747 1027
rect 805 993 811 1053
rect 821 1027 827 1053
rect 805 987 827 993
rect 757 827 763 853
rect 773 833 779 933
rect 821 853 827 987
rect 885 853 891 1253
rect 917 1193 923 1273
rect 933 1247 939 1473
rect 965 1467 971 1613
rect 997 1607 1011 1613
rect 965 1227 971 1273
rect 917 1187 939 1193
rect 933 1027 939 1187
rect 965 1087 971 1133
rect 981 873 987 1593
rect 1005 1493 1011 1607
rect 997 1487 1011 1493
rect 1045 1493 1051 1667
rect 1045 1487 1083 1493
rect 997 1413 1003 1487
rect 1045 1453 1051 1473
rect 1013 1447 1051 1453
rect 997 1407 1019 1413
rect 1013 1293 1019 1407
rect 997 1287 1019 1293
rect 997 1247 1003 1287
rect 1013 1207 1019 1233
rect 997 987 1003 1193
rect 1013 1033 1019 1093
rect 1045 1067 1051 1433
rect 1077 1327 1083 1487
rect 1109 1347 1115 1653
rect 1125 1607 1131 1853
rect 1141 1667 1147 1853
rect 1221 1733 1227 2007
rect 1237 1847 1243 1893
rect 1253 1833 1259 2033
rect 1285 1847 1291 2053
rect 1301 1847 1307 2127
rect 1317 2013 1323 2133
rect 1397 2127 1403 2333
rect 1429 2327 1435 2593
rect 1445 2427 1483 2433
rect 1493 2413 1499 2593
rect 1573 2587 1579 2653
rect 1605 2547 1611 2733
rect 1621 2707 1627 3047
rect 1637 2727 1643 2993
rect 1653 2807 1659 3033
rect 1717 2987 1723 3073
rect 1733 3067 1739 3107
rect 1733 3007 1739 3053
rect 1829 3027 1835 3073
rect 1845 3013 1851 3147
rect 1893 3067 1899 3133
rect 1909 3113 1915 3233
rect 1925 3133 1931 3247
rect 1973 3227 1979 3267
rect 2021 3153 2027 3307
rect 2133 3247 2139 3307
rect 2053 3207 2059 3233
rect 2149 3227 2155 3473
rect 2165 3467 2187 3473
rect 2165 3447 2203 3453
rect 2469 3433 2475 3453
rect 2485 3447 2491 3473
rect 2469 3427 2491 3433
rect 2501 3387 2507 3453
rect 2021 3147 2043 3153
rect 1925 3127 2027 3133
rect 1909 3107 1947 3113
rect 1893 3033 1899 3053
rect 1909 3047 1915 3073
rect 1941 3067 1947 3107
rect 1973 3067 1995 3073
rect 2021 3067 2027 3127
rect 2037 3113 2043 3147
rect 2085 3133 2091 3193
rect 2077 3127 2091 3133
rect 2037 3107 2059 3113
rect 1925 3047 1947 3053
rect 1925 3033 1931 3047
rect 1797 3007 1851 3013
rect 1877 3007 1883 3033
rect 1893 3027 1931 3033
rect 1717 2873 1723 2913
rect 1669 2847 1675 2873
rect 1701 2867 1723 2873
rect 1701 2733 1707 2867
rect 1733 2807 1739 2873
rect 1749 2793 1755 2893
rect 1733 2787 1755 2793
rect 1765 2847 1787 2853
rect 1701 2727 1723 2733
rect 1621 2667 1627 2693
rect 1717 2667 1723 2727
rect 1733 2667 1739 2787
rect 1445 2407 1499 2413
rect 1445 2387 1451 2407
rect 1541 2387 1547 2413
rect 1557 2407 1563 2453
rect 1653 2333 1659 2613
rect 1669 2427 1707 2433
rect 1717 2393 1723 2653
rect 1733 2533 1739 2653
rect 1749 2567 1755 2673
rect 1765 2647 1771 2847
rect 1781 2687 1787 2833
rect 1797 2807 1803 3007
rect 1941 2907 1947 3033
rect 1813 2827 1819 2853
rect 1829 2827 1835 2893
rect 2021 2887 2027 3033
rect 2053 2893 2059 3107
rect 2077 3013 2083 3127
rect 2101 3013 2107 3173
rect 2197 3087 2203 3293
rect 2245 3227 2251 3253
rect 2229 3167 2235 3213
rect 2213 3127 2251 3133
rect 2197 3047 2203 3073
rect 2213 3067 2219 3127
rect 2213 3033 2219 3053
rect 2229 3047 2235 3073
rect 2245 3053 2251 3127
rect 2261 3067 2267 3193
rect 2357 3107 2363 3213
rect 2389 3207 2395 3373
rect 2405 3227 2411 3273
rect 2437 3207 2443 3233
rect 2517 3227 2523 3473
rect 2533 3467 2555 3473
rect 2533 3427 2539 3453
rect 2629 3227 2635 3393
rect 2709 3287 2715 3473
rect 2741 3447 2747 3473
rect 2709 3227 2715 3273
rect 2613 3187 2619 3213
rect 2357 3067 2363 3093
rect 2245 3047 2267 3053
rect 2213 3027 2251 3033
rect 2261 3013 2267 3047
rect 2325 3013 2331 3053
rect 2077 3007 2091 3013
rect 2101 3007 2139 3013
rect 2261 3007 2331 3013
rect 2085 2967 2091 3007
rect 2037 2887 2059 2893
rect 1909 2867 1995 2873
rect 1877 2833 1883 2853
rect 1909 2847 1915 2867
rect 1845 2827 1867 2833
rect 1877 2827 1915 2833
rect 1989 2827 1995 2867
rect 2037 2833 2043 2887
rect 2021 2827 2043 2833
rect 1845 2813 1851 2827
rect 1813 2807 1851 2813
rect 1781 2573 1787 2673
rect 1797 2647 1803 2793
rect 1813 2667 1819 2733
rect 1813 2627 1819 2653
rect 1829 2587 1835 2793
rect 1861 2787 1867 2813
rect 1877 2807 1899 2813
rect 1845 2687 1899 2693
rect 1845 2667 1851 2687
rect 1861 2667 1883 2673
rect 1893 2667 1899 2687
rect 1861 2627 1867 2653
rect 1909 2627 1915 2827
rect 1925 2767 1931 2813
rect 1925 2647 1931 2753
rect 2021 2747 2027 2813
rect 1781 2567 1867 2573
rect 1733 2527 1755 2533
rect 1669 2387 1723 2393
rect 1749 2353 1755 2527
rect 1845 2407 1851 2513
rect 1861 2427 1867 2567
rect 1877 2393 1883 2553
rect 1941 2527 1947 2693
rect 1957 2607 1963 2693
rect 1869 2387 1883 2393
rect 1413 2247 1419 2273
rect 1333 2027 1339 2053
rect 1429 2027 1435 2273
rect 1509 2093 1515 2213
rect 1525 2133 1531 2313
rect 1541 2267 1547 2293
rect 1541 2247 1579 2253
rect 1589 2187 1595 2333
rect 1605 2327 1659 2333
rect 1733 2347 1755 2353
rect 1605 2207 1611 2327
rect 1733 2313 1739 2347
rect 1621 2307 1739 2313
rect 1621 2267 1627 2307
rect 1637 2213 1643 2273
rect 1637 2207 1675 2213
rect 1733 2207 1739 2273
rect 1749 2267 1755 2293
rect 1749 2227 1755 2253
rect 1845 2207 1851 2373
rect 1525 2127 1547 2133
rect 1509 2087 1523 2093
rect 1317 2007 1339 2013
rect 1381 1907 1387 2013
rect 1477 2007 1483 2033
rect 1517 1953 1523 2087
rect 1541 1987 1547 2127
rect 1573 2047 1643 2053
rect 1573 2027 1579 2047
rect 1509 1947 1523 1953
rect 1317 1833 1323 1873
rect 1429 1867 1435 1933
rect 1253 1827 1323 1833
rect 1157 1727 1227 1733
rect 1157 1607 1163 1727
rect 1189 1467 1195 1653
rect 1205 1607 1211 1633
rect 1221 1607 1227 1673
rect 1237 1627 1243 1693
rect 1333 1687 1339 1853
rect 1269 1607 1275 1633
rect 1301 1607 1307 1673
rect 1237 1467 1243 1493
rect 1269 1467 1291 1473
rect 1253 1407 1259 1453
rect 1125 1367 1163 1373
rect 1093 1227 1115 1233
rect 1077 1187 1083 1213
rect 1093 1187 1099 1227
rect 1125 1213 1131 1367
rect 1237 1253 1243 1353
rect 1229 1247 1243 1253
rect 1109 1207 1131 1213
rect 1109 1173 1115 1207
rect 1077 1167 1115 1173
rect 1077 1047 1083 1167
rect 1157 1127 1179 1133
rect 1013 1027 1035 1033
rect 1029 873 1035 1027
rect 1109 1013 1115 1053
rect 1125 1033 1131 1093
rect 1125 1027 1139 1033
rect 1157 1027 1163 1053
rect 1093 1007 1115 1013
rect 1093 913 1099 1007
rect 1093 907 1115 913
rect 981 867 1003 873
rect 1013 867 1035 873
rect 1109 867 1115 907
rect 1133 873 1139 1027
rect 1125 867 1139 873
rect 805 847 827 853
rect 869 847 891 853
rect 933 847 1003 853
rect 773 827 795 833
rect 741 807 763 813
rect 677 727 699 733
rect 677 647 683 727
rect 725 667 747 673
rect 725 647 731 667
rect 677 407 683 593
rect 725 567 731 633
rect 741 427 747 653
rect 757 647 763 693
rect 789 607 795 827
rect 805 787 811 847
rect 869 693 875 847
rect 917 793 923 833
rect 933 827 939 847
rect 949 807 955 833
rect 917 787 987 793
rect 997 773 1003 847
rect 1013 827 1019 867
rect 869 687 891 693
rect 885 653 891 687
rect 901 667 907 773
rect 981 767 1003 773
rect 949 687 955 753
rect 949 653 955 673
rect 981 653 987 767
rect 837 427 843 653
rect 885 647 955 653
rect 965 647 987 653
rect 901 627 907 647
rect 933 567 939 633
rect 1045 627 1051 773
rect 1125 647 1131 867
rect 1141 767 1147 833
rect 1173 787 1179 1127
rect 1189 993 1195 1053
rect 1205 1027 1211 1213
rect 1229 1133 1235 1247
rect 1229 1127 1243 1133
rect 1221 1067 1227 1093
rect 1237 1013 1243 1127
rect 1253 1067 1259 1233
rect 1285 1227 1291 1433
rect 1301 1353 1307 1573
rect 1317 1393 1323 1533
rect 1365 1513 1371 1733
rect 1429 1653 1435 1853
rect 1461 1667 1467 1873
rect 1509 1787 1515 1947
rect 1557 1887 1563 2013
rect 1573 2007 1595 2013
rect 1557 1827 1563 1853
rect 1605 1813 1611 2033
rect 1637 2027 1643 2047
rect 1621 1927 1627 2013
rect 1637 1987 1643 2013
rect 1669 2007 1675 2207
rect 1765 1913 1771 2193
rect 1869 2093 1875 2387
rect 1893 2267 1899 2433
rect 1925 2407 1931 2433
rect 1957 2387 1963 2413
rect 1973 2367 1979 2713
rect 2037 2707 2043 2813
rect 2133 2773 2139 3007
rect 2149 2887 2187 2893
rect 2149 2827 2155 2887
rect 2165 2827 2171 2873
rect 2181 2847 2187 2887
rect 2277 2873 2283 2993
rect 2197 2867 2267 2873
rect 2277 2867 2299 2873
rect 2197 2833 2203 2867
rect 2181 2827 2203 2833
rect 2261 2827 2267 2867
rect 2181 2813 2187 2827
rect 2149 2807 2187 2813
rect 2101 2767 2139 2773
rect 1989 2667 1995 2693
rect 1989 2627 1995 2653
rect 2005 2427 2011 2593
rect 2053 2527 2059 2653
rect 1989 2327 1995 2413
rect 1925 2307 1963 2313
rect 1893 2227 1899 2253
rect 1869 2087 1883 2093
rect 1781 2027 1787 2053
rect 1781 1967 1787 2013
rect 1877 1953 1883 2087
rect 1861 1947 1883 1953
rect 1717 1907 1771 1913
rect 1717 1873 1723 1907
rect 1709 1867 1723 1873
rect 1589 1807 1611 1813
rect 1429 1647 1467 1653
rect 1397 1553 1403 1633
rect 1461 1567 1467 1647
rect 1477 1647 1563 1653
rect 1477 1607 1483 1647
rect 1493 1607 1499 1633
rect 1509 1553 1515 1613
rect 1525 1607 1531 1633
rect 1541 1607 1547 1633
rect 1557 1627 1563 1647
rect 1397 1547 1515 1553
rect 1557 1513 1563 1613
rect 1365 1507 1419 1513
rect 1557 1507 1579 1513
rect 1413 1467 1419 1507
rect 1381 1393 1387 1453
rect 1413 1407 1419 1453
rect 1429 1447 1435 1473
rect 1461 1393 1467 1433
rect 1477 1413 1483 1473
rect 1573 1467 1579 1507
rect 1525 1447 1547 1453
rect 1573 1413 1579 1453
rect 1477 1407 1579 1413
rect 1317 1387 1339 1393
rect 1381 1387 1467 1393
rect 1301 1347 1315 1353
rect 1309 1213 1315 1347
rect 1301 1207 1315 1213
rect 1301 1067 1307 1207
rect 1333 1153 1339 1387
rect 1317 1147 1339 1153
rect 1317 1107 1323 1147
rect 1253 1033 1259 1053
rect 1285 1047 1307 1053
rect 1285 1033 1291 1047
rect 1253 1027 1291 1033
rect 1301 1013 1307 1033
rect 1237 1007 1307 1013
rect 1189 987 1211 993
rect 1301 987 1307 1007
rect 1205 873 1211 987
rect 1189 867 1211 873
rect 1189 827 1195 867
rect 1237 847 1291 853
rect 1285 813 1291 847
rect 1317 827 1323 1073
rect 1333 1027 1355 1033
rect 1333 813 1339 833
rect 1285 807 1339 813
rect 1173 673 1179 713
rect 1141 667 1179 673
rect 1141 607 1147 667
rect 1189 653 1195 753
rect 1349 673 1355 813
rect 1189 647 1227 653
rect 1157 627 1227 633
rect 1173 333 1179 433
rect 1237 427 1243 673
rect 1301 667 1355 673
rect 1301 433 1307 667
rect 1365 647 1371 793
rect 1381 707 1387 1333
rect 1413 1267 1499 1273
rect 1413 1027 1419 1267
rect 1493 1227 1499 1267
rect 1429 1167 1435 1213
rect 1525 1153 1531 1213
rect 1541 1167 1547 1407
rect 1589 1227 1595 1807
rect 1605 1653 1611 1693
rect 1685 1653 1691 1853
rect 1709 1693 1715 1867
rect 1709 1687 1723 1693
rect 1605 1647 1627 1653
rect 1685 1647 1707 1653
rect 1621 1533 1627 1647
rect 1605 1527 1627 1533
rect 1605 1413 1611 1527
rect 1685 1507 1691 1613
rect 1701 1467 1707 1647
rect 1717 1593 1723 1687
rect 1733 1627 1739 1853
rect 1749 1827 1755 1873
rect 1765 1807 1771 1853
rect 1765 1627 1771 1693
rect 1717 1587 1731 1593
rect 1725 1453 1731 1587
rect 1749 1567 1755 1613
rect 1781 1607 1787 1873
rect 1797 1847 1803 1933
rect 1813 1833 1819 1873
rect 1861 1833 1867 1947
rect 1893 1853 1899 2213
rect 1909 1967 1915 2293
rect 1925 2193 1931 2307
rect 1957 2267 1963 2307
rect 1925 2187 1939 2193
rect 1933 2073 1939 2187
rect 1933 2067 1947 2073
rect 1925 2027 1931 2053
rect 1941 1993 1947 2067
rect 1957 2007 1963 2253
rect 2021 2213 2027 2253
rect 2037 2247 2043 2433
rect 2085 2247 2091 2753
rect 2197 2733 2203 2813
rect 2197 2727 2219 2733
rect 2101 2573 2107 2693
rect 2197 2667 2203 2713
rect 2213 2633 2219 2727
rect 2293 2713 2299 2867
rect 2309 2807 2315 2973
rect 2373 2873 2379 3073
rect 2469 3047 2475 3073
rect 2485 3067 2507 3073
rect 2485 2927 2491 3067
rect 2517 2933 2523 3073
rect 2533 3013 2539 3053
rect 2597 3013 2603 3053
rect 2533 3007 2603 3013
rect 2517 2927 2539 2933
rect 2629 2927 2635 3093
rect 2645 3047 2651 3133
rect 2741 3113 2747 3213
rect 2773 3207 2779 3233
rect 2821 3227 2827 3473
rect 2853 3467 2859 3493
rect 2837 3447 2875 3453
rect 2901 3327 2907 3473
rect 3077 3447 3083 3473
rect 3109 3313 3115 3473
rect 3141 3467 3147 3493
rect 3125 3447 3163 3453
rect 3173 3353 3179 3453
rect 3173 3347 3195 3353
rect 3093 3307 3115 3313
rect 2933 3227 2939 3293
rect 2997 3133 3003 3233
rect 3093 3227 3099 3307
rect 3157 3227 3163 3333
rect 3189 3213 3195 3347
rect 2981 3127 3003 3133
rect 3173 3207 3195 3213
rect 2693 3107 2747 3113
rect 2661 3047 2667 3073
rect 2693 3053 2699 3107
rect 2709 3067 2715 3093
rect 2677 3047 2699 3053
rect 2677 3007 2683 3047
rect 2693 3013 2699 3033
rect 2773 3013 2779 3053
rect 2693 3007 2779 3013
rect 2805 2993 2811 3113
rect 2917 3087 2939 3093
rect 2797 2987 2811 2993
rect 2373 2867 2427 2873
rect 2341 2847 2379 2853
rect 2341 2827 2347 2847
rect 2373 2827 2379 2847
rect 2261 2707 2299 2713
rect 2205 2627 2219 2633
rect 2117 2573 2123 2593
rect 2101 2567 2123 2573
rect 2101 2373 2107 2413
rect 2117 2407 2123 2567
rect 2205 2493 2211 2627
rect 2205 2487 2219 2493
rect 2229 2487 2235 2673
rect 2245 2573 2251 2673
rect 2261 2667 2267 2707
rect 2357 2667 2363 2733
rect 2405 2713 2411 2813
rect 2421 2807 2427 2867
rect 2469 2827 2491 2833
rect 2517 2807 2523 2873
rect 2405 2707 2475 2713
rect 2261 2613 2267 2653
rect 2325 2613 2331 2653
rect 2261 2607 2331 2613
rect 2373 2607 2379 2673
rect 2245 2567 2259 2573
rect 2213 2433 2219 2487
rect 2253 2453 2259 2567
rect 2277 2467 2347 2473
rect 2253 2447 2267 2453
rect 2213 2427 2235 2433
rect 2101 2367 2171 2373
rect 2133 2273 2139 2353
rect 2117 2267 2139 2273
rect 2165 2267 2171 2367
rect 2213 2287 2219 2413
rect 2117 2247 2123 2267
rect 2005 2027 2011 2213
rect 2021 2207 2043 2213
rect 2133 2207 2139 2253
rect 2037 2073 2043 2207
rect 2229 2187 2235 2427
rect 2245 2327 2251 2413
rect 2261 2407 2267 2447
rect 2277 2427 2283 2467
rect 2341 2427 2347 2467
rect 2373 2407 2395 2413
rect 2373 2387 2395 2393
rect 2021 2067 2043 2073
rect 2021 2007 2027 2067
rect 1925 1867 1931 1993
rect 1941 1987 1979 1993
rect 1973 1867 1979 1987
rect 2037 1873 2043 2033
rect 2053 1927 2059 2013
rect 2069 1887 2075 2013
rect 2085 2007 2091 2033
rect 2101 2007 2107 2053
rect 2117 1973 2123 2033
rect 2213 2027 2219 2053
rect 2109 1967 2123 1973
rect 2037 1867 2075 1873
rect 1893 1847 1915 1853
rect 1813 1827 1835 1833
rect 1861 1827 1883 1833
rect 1829 1733 1835 1827
rect 1813 1727 1835 1733
rect 1813 1553 1819 1727
rect 1877 1687 1883 1827
rect 1909 1653 1915 1847
rect 2053 1813 2059 1853
rect 2045 1807 2059 1813
rect 1893 1647 1915 1653
rect 1861 1567 1867 1633
rect 1717 1447 1731 1453
rect 1749 1547 1819 1553
rect 1893 1553 1899 1647
rect 1941 1593 1947 1693
rect 1957 1647 1995 1653
rect 1957 1627 1963 1647
rect 1941 1587 1955 1593
rect 1893 1547 1915 1553
rect 1717 1413 1723 1447
rect 1605 1407 1643 1413
rect 1573 1153 1579 1213
rect 1525 1147 1579 1153
rect 1445 1033 1451 1113
rect 1509 1067 1515 1113
rect 1461 1047 1515 1053
rect 1445 1027 1467 1033
rect 1477 1027 1499 1033
rect 1445 773 1451 993
rect 1461 827 1467 1027
rect 1509 1013 1515 1047
rect 1573 1013 1579 1053
rect 1477 987 1483 1013
rect 1509 1007 1579 1013
rect 1605 993 1611 1053
rect 1597 987 1611 993
rect 1597 873 1603 987
rect 1557 867 1603 873
rect 1557 807 1563 867
rect 1413 767 1451 773
rect 1605 767 1611 853
rect 1301 427 1339 433
rect 1381 407 1387 673
rect 1413 627 1419 767
rect 1621 727 1627 1173
rect 1637 827 1643 1407
rect 1685 1407 1723 1413
rect 1653 1033 1659 1253
rect 1685 1187 1691 1407
rect 1749 1313 1755 1547
rect 1813 1467 1819 1533
rect 1909 1467 1915 1547
rect 1765 1447 1819 1453
rect 1781 1407 1787 1433
rect 1797 1367 1803 1433
rect 1813 1413 1819 1447
rect 1877 1413 1883 1453
rect 1925 1447 1931 1493
rect 1949 1433 1955 1587
rect 1973 1507 1979 1633
rect 1989 1627 1995 1647
rect 1989 1587 1995 1613
rect 2021 1607 2027 1693
rect 2045 1673 2051 1807
rect 2045 1667 2059 1673
rect 2037 1587 2043 1633
rect 2053 1607 2059 1667
rect 2069 1627 2075 1867
rect 2109 1793 2115 1967
rect 2133 1927 2139 2013
rect 2149 1913 2155 1973
rect 2133 1907 2155 1913
rect 2133 1813 2139 1907
rect 2165 1867 2171 2013
rect 2245 1967 2251 2253
rect 2325 2213 2331 2293
rect 2325 2207 2347 2213
rect 2325 2027 2331 2193
rect 2357 2167 2363 2253
rect 2357 2007 2363 2033
rect 2373 2007 2379 2387
rect 2405 2373 2411 2653
rect 2437 2627 2443 2653
rect 2469 2647 2475 2707
rect 2485 2687 2491 2773
rect 2501 2667 2507 2693
rect 2517 2633 2523 2713
rect 2533 2667 2539 2927
rect 2797 2873 2803 2987
rect 2821 2967 2827 3073
rect 2869 3047 2891 3053
rect 2757 2867 2803 2873
rect 2645 2827 2651 2853
rect 2629 2687 2635 2813
rect 2645 2787 2651 2813
rect 2741 2707 2747 2813
rect 2757 2693 2763 2867
rect 2789 2827 2795 2853
rect 2773 2747 2779 2813
rect 2821 2707 2827 2953
rect 2917 2873 2923 3073
rect 2933 3067 2939 3087
rect 2901 2867 2923 2873
rect 2741 2687 2763 2693
rect 2501 2627 2523 2633
rect 2405 2367 2475 2373
rect 2437 2207 2443 2253
rect 2469 2073 2475 2367
rect 2501 2347 2507 2627
rect 2533 2613 2539 2653
rect 2597 2613 2603 2653
rect 2533 2607 2603 2613
rect 2533 2407 2539 2573
rect 2629 2493 2635 2673
rect 2645 2587 2651 2673
rect 2629 2487 2683 2493
rect 2565 2467 2635 2473
rect 2565 2427 2571 2467
rect 2629 2427 2635 2467
rect 2549 2313 2555 2413
rect 2565 2373 2571 2413
rect 2677 2393 2683 2487
rect 2693 2407 2699 2653
rect 2661 2387 2683 2393
rect 2565 2367 2619 2373
rect 2517 2307 2555 2313
rect 2517 2213 2523 2307
rect 2517 2207 2539 2213
rect 2389 2067 2475 2073
rect 2389 1873 2395 2067
rect 2485 1967 2491 2013
rect 2517 2007 2523 2073
rect 2533 2007 2539 2207
rect 2581 2167 2587 2253
rect 2613 2087 2619 2367
rect 2629 2267 2635 2313
rect 2661 2253 2667 2387
rect 2645 2247 2667 2253
rect 2549 2067 2619 2073
rect 2549 2027 2555 2067
rect 2613 2027 2619 2067
rect 2261 1833 2267 1853
rect 2277 1847 2283 1873
rect 2293 1833 2299 1873
rect 2373 1867 2395 1873
rect 2261 1827 2299 1833
rect 2133 1807 2155 1813
rect 2109 1787 2123 1793
rect 2085 1607 2091 1633
rect 2101 1627 2107 1693
rect 2117 1627 2123 1787
rect 2149 1673 2155 1807
rect 2325 1793 2331 1833
rect 2133 1667 2155 1673
rect 2317 1787 2331 1793
rect 2133 1613 2139 1667
rect 2213 1647 2299 1653
rect 2101 1607 2139 1613
rect 2101 1513 2107 1607
rect 2181 1587 2187 1633
rect 2213 1607 2219 1647
rect 2245 1627 2267 1633
rect 2293 1627 2299 1647
rect 2101 1507 2123 1513
rect 1813 1407 1883 1413
rect 1941 1427 1955 1433
rect 1749 1307 1803 1313
rect 1669 1067 1675 1113
rect 1653 1027 1667 1033
rect 1661 893 1667 1027
rect 1653 887 1667 893
rect 1653 847 1659 887
rect 1445 667 1451 713
rect 1637 667 1643 713
rect 1685 673 1691 1153
rect 1701 1027 1707 1073
rect 1717 1047 1723 1233
rect 1733 1207 1739 1273
rect 1749 1227 1755 1253
rect 1733 827 1739 1073
rect 1765 1067 1771 1213
rect 1797 1147 1803 1307
rect 1845 1227 1851 1273
rect 1941 1233 1947 1427
rect 1973 1367 1979 1473
rect 2021 1467 2027 1493
rect 2117 1467 2123 1507
rect 2005 1413 2011 1433
rect 2085 1413 2091 1453
rect 2005 1407 2091 1413
rect 1973 1267 2059 1273
rect 1925 1227 1947 1233
rect 1925 1153 1931 1227
rect 1861 1147 1931 1153
rect 1781 1073 1787 1113
rect 1861 1073 1867 1147
rect 1781 1067 1867 1073
rect 1749 947 1755 1053
rect 1781 1027 1787 1053
rect 1845 827 1851 1067
rect 1893 1047 1899 1093
rect 1925 1067 1931 1133
rect 1941 893 1947 1213
rect 1957 1187 1963 1233
rect 1973 1173 1979 1267
rect 1989 1227 1995 1253
rect 2053 1227 2059 1267
rect 2133 1253 2139 1473
rect 2229 1467 2235 1573
rect 2245 1533 2251 1613
rect 2261 1607 2283 1613
rect 2293 1567 2299 1613
rect 2317 1573 2323 1787
rect 2341 1613 2347 1853
rect 2357 1627 2363 1733
rect 2341 1607 2363 1613
rect 2317 1567 2331 1573
rect 2245 1527 2315 1533
rect 2197 1367 2203 1453
rect 2261 1353 2267 1473
rect 2309 1447 2315 1527
rect 2181 1347 2267 1353
rect 2101 1247 2139 1253
rect 2085 1193 2091 1213
rect 2101 1207 2107 1247
rect 2117 1193 2123 1213
rect 2133 1193 2139 1213
rect 2085 1187 2139 1193
rect 1973 1167 2027 1173
rect 1957 987 1963 1073
rect 1989 1047 1995 1093
rect 2021 1047 2027 1167
rect 1941 887 1963 893
rect 1685 667 1723 673
rect 1813 667 1819 693
rect 1893 673 1899 813
rect 1957 793 1963 887
rect 1941 787 1963 793
rect 1941 673 1947 787
rect 1861 667 1899 673
rect 1909 667 1947 673
rect 1445 427 1483 433
rect 1509 427 1515 653
rect 1605 627 1611 653
rect 1685 513 1691 653
rect 1637 507 1691 513
rect 1477 413 1483 427
rect 1477 407 1547 413
rect 1157 327 1179 333
rect 1157 267 1163 327
rect 1493 313 1499 393
rect 1493 307 1531 313
rect 1333 267 1339 293
rect 1253 173 1259 253
rect 1317 227 1323 253
rect 1333 173 1339 253
rect 1477 247 1483 273
rect 1493 233 1499 307
rect 1477 227 1499 233
rect 1509 227 1515 293
rect 1525 267 1531 307
rect 1589 293 1595 433
rect 1637 427 1643 507
rect 1717 447 1723 667
rect 1669 367 1675 413
rect 1557 287 1595 293
rect 1589 267 1595 287
rect 1717 273 1723 433
rect 1829 407 1835 433
rect 1861 367 1867 667
rect 1877 613 1883 653
rect 1893 627 1899 653
rect 1909 613 1915 667
rect 1877 607 1915 613
rect 1925 407 1931 653
rect 1957 647 1963 733
rect 1989 647 1995 833
rect 2037 813 2043 1053
rect 2085 1047 2107 1053
rect 2149 1013 2155 1253
rect 2181 1213 2187 1347
rect 2261 1313 2267 1333
rect 2213 1307 2267 1313
rect 2213 1227 2219 1307
rect 2181 1207 2203 1213
rect 2197 1147 2203 1207
rect 2181 1067 2203 1073
rect 2229 1047 2235 1233
rect 2245 1207 2251 1293
rect 2261 1227 2267 1307
rect 2245 1027 2251 1073
rect 2277 1067 2283 1213
rect 2293 1207 2299 1233
rect 2309 1207 2315 1253
rect 2325 1053 2331 1567
rect 2341 1327 2347 1593
rect 2357 1207 2363 1607
rect 2373 1593 2379 1867
rect 2405 1853 2411 1933
rect 2645 1927 2651 2247
rect 2693 2213 2699 2393
rect 2725 2387 2731 2413
rect 2741 2313 2747 2687
rect 2773 2507 2779 2673
rect 2789 2607 2795 2673
rect 2805 2613 2811 2653
rect 2869 2613 2875 2653
rect 2805 2607 2875 2613
rect 2773 2467 2843 2473
rect 2773 2427 2779 2467
rect 2837 2427 2843 2467
rect 2757 2367 2763 2413
rect 2741 2307 2811 2313
rect 2773 2213 2779 2253
rect 2693 2207 2779 2213
rect 2677 2007 2683 2193
rect 2805 2113 2811 2307
rect 2869 2273 2875 2313
rect 2901 2293 2907 2867
rect 2917 2827 2923 2853
rect 2949 2787 2955 3053
rect 2981 2993 2987 3127
rect 3077 3047 3083 3113
rect 3141 3047 3147 3093
rect 3157 3007 3163 3053
rect 2965 2987 2987 2993
rect 2965 2947 2971 2987
rect 2933 2667 2939 2713
rect 2965 2693 2971 2933
rect 2981 2813 2987 2973
rect 3013 2827 3019 2893
rect 2981 2807 3003 2813
rect 2965 2687 2987 2693
rect 2965 2427 2971 2593
rect 2853 2267 2875 2273
rect 2893 2287 2907 2293
rect 2853 2153 2859 2267
rect 2893 2173 2899 2287
rect 2949 2273 2955 2413
rect 2981 2407 2987 2687
rect 3029 2673 3035 2813
rect 3061 2807 3067 2853
rect 3077 2827 3115 2833
rect 3173 2813 3179 3207
rect 3189 3073 3195 3113
rect 3237 3073 3243 3493
rect 3189 3067 3211 3073
rect 3237 3067 3275 3073
rect 3221 3047 3259 3053
rect 3005 2667 3035 2673
rect 3005 2453 3011 2667
rect 2997 2447 3011 2453
rect 2997 2407 3003 2447
rect 3029 2407 3035 2653
rect 3045 2427 3083 2433
rect 3093 2413 3099 2813
rect 3157 2807 3179 2813
rect 3157 2767 3163 2807
rect 3125 2587 3131 2653
rect 3061 2407 3099 2413
rect 2917 2267 2955 2273
rect 2917 2193 2923 2267
rect 2949 2233 2955 2253
rect 2965 2247 2971 2373
rect 3061 2313 3067 2407
rect 3029 2307 3067 2313
rect 2981 2267 2987 2293
rect 2997 2233 3003 2253
rect 2949 2227 3003 2233
rect 2917 2187 2939 2193
rect 2893 2167 2907 2173
rect 2853 2147 2875 2153
rect 2805 2107 2827 2113
rect 2421 1907 2523 1913
rect 2421 1867 2427 1907
rect 2453 1867 2459 1893
rect 2389 1607 2395 1853
rect 2405 1847 2427 1853
rect 2373 1587 2395 1593
rect 2389 1453 2395 1587
rect 2389 1447 2411 1453
rect 2421 1447 2427 1847
rect 2469 1827 2475 1853
rect 2485 1653 2491 1873
rect 2501 1827 2507 1853
rect 2517 1813 2523 1907
rect 2517 1807 2539 1813
rect 2533 1693 2539 1807
rect 2613 1713 2619 1873
rect 2661 1847 2667 1893
rect 2741 1753 2747 2093
rect 2773 2027 2779 2053
rect 2821 2013 2827 2107
rect 2869 2027 2875 2147
rect 2805 2007 2827 2013
rect 2581 1707 2619 1713
rect 2725 1747 2747 1753
rect 2533 1687 2555 1693
rect 2469 1627 2475 1653
rect 2485 1647 2539 1653
rect 2501 1627 2523 1633
rect 2469 1547 2475 1613
rect 2501 1587 2507 1613
rect 2533 1607 2539 1647
rect 2549 1593 2555 1687
rect 2581 1607 2587 1707
rect 2533 1587 2555 1593
rect 2629 1587 2635 1633
rect 2725 1613 2731 1747
rect 2757 1627 2763 1993
rect 2805 1853 2811 2007
rect 2901 1987 2907 2167
rect 2933 2053 2939 2187
rect 2917 2047 2939 2053
rect 2773 1847 2811 1853
rect 2773 1827 2779 1847
rect 2821 1673 2827 1873
rect 2837 1847 2843 1973
rect 2917 1847 2923 2047
rect 2965 2007 2971 2053
rect 2981 2027 3019 2033
rect 3029 2013 3035 2307
rect 3077 2027 3083 2273
rect 3125 2247 3131 2293
rect 3157 2187 3163 2713
rect 3221 2607 3227 2833
rect 3269 2787 3275 3067
rect 3301 2827 3339 2833
rect 3285 2733 3291 2813
rect 3317 2787 3323 2813
rect 3253 2727 3291 2733
rect 3253 2647 3259 2727
rect 3349 2607 3355 2653
rect 3269 2247 3275 2373
rect 2997 2007 3035 2013
rect 3205 2007 3243 2013
rect 2997 1967 3003 2007
rect 3205 1887 3259 1893
rect 2805 1667 2827 1673
rect 2725 1607 2747 1613
rect 2357 1067 2363 1153
rect 2405 1067 2411 1447
rect 2437 1313 2443 1493
rect 2533 1467 2539 1587
rect 2565 1427 2571 1473
rect 2437 1307 2451 1313
rect 2421 1227 2427 1293
rect 2445 1213 2451 1307
rect 2581 1287 2587 1473
rect 2693 1467 2699 1553
rect 2597 1413 2603 1453
rect 2661 1413 2667 1453
rect 2597 1407 2667 1413
rect 2645 1307 2731 1313
rect 2517 1227 2523 1253
rect 2437 1207 2451 1213
rect 2261 1047 2331 1053
rect 2101 1007 2155 1013
rect 2053 827 2059 853
rect 2037 807 2075 813
rect 2101 767 2107 1007
rect 2133 813 2139 853
rect 2149 827 2155 933
rect 2261 927 2267 1047
rect 2421 1027 2427 1053
rect 2277 907 2363 913
rect 2277 827 2283 907
rect 2133 807 2155 813
rect 2053 687 2123 693
rect 2053 667 2059 687
rect 2069 667 2091 673
rect 1957 427 1963 453
rect 2021 427 2027 633
rect 2037 427 2043 453
rect 2085 427 2091 653
rect 2117 647 2123 687
rect 2133 667 2139 693
rect 2149 647 2155 807
rect 2181 787 2187 813
rect 2341 807 2347 833
rect 2357 827 2363 907
rect 2437 893 2443 1207
rect 2517 1047 2523 1073
rect 2421 887 2443 893
rect 2357 793 2363 813
rect 2421 807 2427 887
rect 2437 847 2491 853
rect 2437 827 2443 847
rect 2469 793 2475 833
rect 2357 787 2475 793
rect 2421 753 2427 773
rect 2437 753 2443 773
rect 2421 747 2443 753
rect 2373 727 2427 733
rect 2229 667 2235 713
rect 2373 653 2379 727
rect 2389 667 2395 713
rect 2421 667 2427 727
rect 2437 667 2443 747
rect 2165 627 2171 653
rect 2277 427 2283 653
rect 2341 613 2347 653
rect 2373 647 2395 653
rect 2405 613 2411 653
rect 2485 647 2491 847
rect 2501 787 2507 813
rect 2517 687 2523 873
rect 2549 747 2555 1233
rect 2645 1227 2651 1307
rect 2709 1233 2715 1293
rect 2693 1227 2715 1233
rect 2725 1227 2731 1307
rect 2741 1247 2747 1607
rect 2773 1547 2779 1633
rect 2805 1573 2811 1667
rect 3013 1653 3019 1873
rect 2949 1627 2955 1653
rect 2997 1647 3019 1653
rect 2805 1567 2827 1573
rect 2581 1027 2587 1053
rect 2597 767 2603 1213
rect 2693 1153 2699 1227
rect 2645 1147 2699 1153
rect 2613 1047 2619 1093
rect 2629 867 2635 1073
rect 2645 1047 2651 1147
rect 2725 1087 2731 1213
rect 2661 1067 2699 1073
rect 2661 1027 2667 1053
rect 2613 693 2619 833
rect 2629 827 2683 833
rect 2677 727 2683 827
rect 2693 807 2699 1067
rect 2773 1013 2779 1533
rect 2821 1207 2827 1567
rect 2853 1527 2859 1613
rect 2933 1467 2939 1613
rect 2997 1527 3003 1647
rect 3013 1627 3067 1633
rect 3077 1627 3083 1653
rect 3109 1633 3115 1853
rect 3109 1627 3147 1633
rect 3013 1587 3035 1593
rect 3045 1573 3051 1613
rect 3061 1593 3067 1627
rect 3061 1587 3099 1593
rect 3029 1567 3051 1573
rect 3029 1467 3035 1567
rect 3093 1547 3099 1587
rect 3109 1553 3115 1613
rect 3173 1607 3179 1853
rect 3205 1607 3211 1887
rect 3237 1867 3259 1873
rect 3109 1547 3131 1553
rect 3157 1547 3163 1593
rect 3061 1467 3067 1533
rect 2837 1267 2939 1273
rect 2837 1207 2843 1267
rect 2853 1047 2859 1233
rect 2869 1207 2875 1253
rect 2885 1207 2891 1233
rect 2933 1227 2939 1267
rect 2981 1207 2987 1453
rect 3125 1393 3131 1547
rect 3109 1387 3131 1393
rect 3045 1227 3067 1233
rect 2997 1107 3003 1213
rect 2901 1047 2939 1053
rect 2725 1007 2779 1013
rect 2725 747 2731 1007
rect 2821 807 2827 833
rect 2597 687 2619 693
rect 2597 673 2603 687
rect 2341 607 2411 613
rect 2501 607 2507 673
rect 2549 667 2603 673
rect 2549 627 2555 667
rect 2341 433 2347 607
rect 2373 467 2443 473
rect 2021 407 2043 413
rect 2181 387 2187 413
rect 1717 267 1739 273
rect 1589 227 1595 253
rect 1733 247 1739 267
rect 1749 247 1755 273
rect 2293 267 2299 433
rect 2341 427 2363 433
rect 2373 427 2379 467
rect 2437 427 2443 467
rect 2533 427 2539 453
rect 2565 427 2571 653
rect 2613 607 2619 673
rect 2341 387 2347 413
rect 2357 407 2363 427
rect 2613 393 2619 593
rect 2629 567 2635 673
rect 2645 613 2651 653
rect 2709 613 2715 653
rect 2645 607 2715 613
rect 2629 427 2699 433
rect 2629 407 2635 427
rect 2661 393 2667 413
rect 2501 267 2507 393
rect 2613 387 2667 393
rect 2533 267 2539 353
rect 2693 267 2699 427
rect 2741 407 2747 633
rect 2757 587 2763 673
rect 2837 667 2843 693
rect 2853 667 2859 873
rect 2885 693 2891 833
rect 2901 727 2907 1047
rect 2965 933 2971 1093
rect 3061 1027 3067 1053
rect 3109 1033 3115 1387
rect 3157 1227 3163 1453
rect 3221 1447 3227 1493
rect 3237 1227 3243 1867
rect 3253 1847 3291 1853
rect 3301 1827 3307 1873
rect 3397 1867 3403 1893
rect 3365 1807 3371 1853
rect 3365 1627 3371 1653
rect 3397 1627 3403 1853
rect 3429 1827 3435 1853
rect 3477 1807 3483 1853
rect 3493 1673 3499 1873
rect 3461 1667 3499 1673
rect 3429 1613 3435 1633
rect 3285 1453 3291 1613
rect 3397 1607 3435 1613
rect 3397 1547 3403 1607
rect 3461 1573 3467 1667
rect 3477 1627 3483 1653
rect 3429 1567 3467 1573
rect 3349 1487 3387 1493
rect 3349 1467 3355 1487
rect 3381 1473 3387 1487
rect 3365 1453 3371 1473
rect 3381 1467 3403 1473
rect 3285 1447 3371 1453
rect 3429 1247 3435 1567
rect 3477 1253 3483 1613
rect 3509 1413 3515 1453
rect 3509 1407 3531 1413
rect 3525 1293 3531 1407
rect 3509 1287 3531 1293
rect 3253 1227 3307 1233
rect 3125 1047 3131 1213
rect 3253 1187 3259 1227
rect 3141 1033 3147 1093
rect 3109 1027 3147 1033
rect 2965 927 2987 933
rect 2917 807 2923 873
rect 2949 807 2955 833
rect 2981 733 2987 927
rect 3109 867 3115 1027
rect 3157 973 3163 1113
rect 3317 1053 3323 1213
rect 3365 1133 3371 1213
rect 3381 1167 3387 1233
rect 3445 1227 3451 1253
rect 3461 1247 3483 1253
rect 3461 1213 3467 1247
rect 3413 1153 3419 1213
rect 3445 1207 3467 1213
rect 3445 1167 3451 1207
rect 3477 1153 3483 1233
rect 3493 1227 3499 1253
rect 3413 1147 3483 1153
rect 3509 1153 3515 1287
rect 3573 1267 3643 1273
rect 3541 1167 3547 1213
rect 3557 1207 3563 1253
rect 3573 1227 3579 1267
rect 3637 1227 3643 1267
rect 3669 1187 3675 1213
rect 3509 1147 3611 1153
rect 3365 1127 3387 1133
rect 3333 1107 3371 1113
rect 3333 1067 3339 1107
rect 3189 1027 3195 1053
rect 3141 967 3163 973
rect 3077 827 3083 853
rect 3141 827 3147 967
rect 3173 807 3179 873
rect 3205 827 3211 853
rect 3269 827 3275 1053
rect 3285 1027 3291 1053
rect 3317 1047 3339 1053
rect 3365 1013 3371 1107
rect 3381 1073 3387 1127
rect 3381 1067 3403 1073
rect 3413 1053 3419 1147
rect 3509 1093 3515 1147
rect 3461 1087 3515 1093
rect 3381 1027 3387 1053
rect 3397 1047 3419 1053
rect 3461 1047 3499 1053
rect 3349 1007 3371 1013
rect 3285 833 3291 893
rect 3349 873 3355 1007
rect 3349 867 3371 873
rect 3285 827 3339 833
rect 2965 727 2987 733
rect 2869 687 2891 693
rect 2869 653 2875 687
rect 2965 667 2971 727
rect 3157 673 3163 793
rect 3125 667 3163 673
rect 2773 427 2779 653
rect 2789 647 2875 653
rect 2933 573 2939 653
rect 3013 573 3019 653
rect 3125 647 3131 667
rect 3157 653 3163 667
rect 2933 567 3019 573
rect 2917 467 2987 473
rect 2805 447 2891 453
rect 2821 393 2827 433
rect 2837 427 2859 433
rect 2853 393 2859 427
rect 2885 407 2891 447
rect 2917 427 2923 467
rect 2981 427 2987 467
rect 3141 433 3147 653
rect 3157 647 3211 653
rect 3221 613 3227 673
rect 3205 607 3227 613
rect 3237 667 3323 673
rect 3205 433 3211 607
rect 3237 447 3243 667
rect 3333 653 3339 673
rect 3349 667 3355 813
rect 3365 807 3371 867
rect 3381 813 3387 833
rect 3397 827 3403 1047
rect 3509 827 3515 1087
rect 3605 1067 3611 1147
rect 3557 833 3563 1053
rect 3541 827 3563 833
rect 3605 827 3611 1053
rect 3381 807 3467 813
rect 2901 393 2907 413
rect 2821 387 2843 393
rect 2853 387 2907 393
rect 3013 387 3019 433
rect 3077 427 3115 433
rect 3141 427 3163 433
rect 3205 427 3227 433
rect 3253 427 3259 653
rect 3269 647 3339 653
rect 3269 427 3275 453
rect 3301 433 3307 633
rect 3333 627 3339 647
rect 3349 613 3355 653
rect 3413 613 3419 653
rect 3461 633 3467 807
rect 3541 733 3547 827
rect 3541 727 3563 733
rect 3349 607 3419 613
rect 3445 627 3467 633
rect 3317 467 3355 473
rect 3317 433 3323 467
rect 3301 427 3323 433
rect 3333 427 3339 453
rect 3045 393 3051 413
rect 3077 407 3083 427
rect 3109 393 3115 413
rect 3045 387 3115 393
rect 2725 267 2731 293
rect 2629 187 2635 253
rect 2645 227 2651 253
rect 2725 213 2731 253
rect 2789 213 2795 253
rect 2821 227 2827 273
rect 2725 207 2795 213
rect 2837 187 2843 387
rect 2869 247 2875 293
rect 2917 267 2923 353
rect 2949 267 2955 373
rect 2965 247 2971 293
rect 2981 227 2987 293
rect 3045 267 3051 387
rect 3157 327 3163 413
rect 3221 387 3227 427
rect 3061 247 3067 293
rect 3221 267 3227 373
rect 3317 367 3323 413
rect 3349 407 3355 467
rect 3381 427 3387 493
rect 3445 387 3451 627
rect 3493 407 3499 433
rect 3509 407 3515 653
rect 3525 647 3531 693
rect 3557 627 3563 727
rect 3573 667 3579 813
rect 3573 487 3579 653
rect 3589 627 3595 653
rect 3525 467 3595 473
rect 3525 427 3531 467
rect 3589 427 3595 467
rect 3621 387 3627 413
rect 3077 227 3083 253
rect 1253 167 1339 173
rect 3708 74 3748 3606
rect 3756 26 3796 3654
<< metal3 >>
rect 1475 3565 1645 3575
rect 1795 3505 2125 3515
rect 819 3485 1581 3495
rect 1603 3485 1757 3495
rect 1571 3475 1581 3485
rect 1795 3475 1805 3505
rect 1571 3465 1805 3475
rect 2115 3475 2125 3505
rect 2595 3505 2813 3515
rect 2211 3485 2493 3495
rect 2211 3475 2221 3485
rect 2115 3465 2221 3475
rect 2483 3475 2493 3485
rect 2595 3475 2605 3505
rect 2803 3495 2813 3505
rect 2803 3485 3245 3495
rect 2483 3465 2605 3475
rect 1139 3445 1197 3455
rect 1827 3445 2093 3455
rect 1187 3435 1197 3445
rect 1555 3435 1837 3445
rect 2083 3435 2093 3445
rect 2243 3445 2797 3455
rect 2243 3435 2253 3445
rect 2787 3435 2797 3445
rect 3027 3445 3181 3455
rect 3027 3435 3037 3445
rect 1187 3425 1565 3435
rect 2083 3425 2253 3435
rect 2483 3425 2541 3435
rect 2787 3425 3037 3435
rect 1603 3405 1949 3415
rect 1987 3385 2349 3395
rect 2499 3385 2637 3395
rect 1987 3375 1997 3385
rect 1475 3365 1997 3375
rect 2339 3375 2349 3385
rect 2339 3365 2397 3375
rect 2675 3345 2861 3355
rect 1827 3335 2045 3345
rect 2675 3335 2685 3345
rect 1715 3325 1837 3335
rect 2035 3325 2685 3335
rect 2851 3335 2861 3345
rect 2851 3325 3165 3335
rect 1859 3305 2013 3315
rect 739 3285 1293 3295
rect 2195 3285 2941 3295
rect 739 3275 749 3285
rect 691 3265 749 3275
rect 1283 3275 1293 3285
rect 1283 3265 1533 3275
rect 2403 3265 2461 3275
rect 2659 3265 2717 3275
rect 2451 3255 2669 3265
rect 403 3245 621 3255
rect 1667 3245 1805 3255
rect 1843 3245 1917 3255
rect 2131 3245 2253 3255
rect 1667 3235 1677 3245
rect 707 3225 925 3235
rect 1043 3225 1261 3235
rect 1443 3225 1677 3235
rect 1795 3235 1805 3245
rect 1795 3225 3005 3235
rect 1443 3195 1453 3225
rect 547 3185 685 3195
rect 851 3185 989 3195
rect 1027 3185 1453 3195
rect 1699 3185 1885 3195
rect 2083 3185 2621 3195
rect 1027 3175 1037 3185
rect 835 3165 1037 3175
rect 2099 3165 2237 3175
rect 803 3145 1117 3155
rect 1235 3145 1469 3155
rect 1731 3145 1917 3155
rect 2323 3145 2605 3155
rect 2323 3135 2333 3145
rect 1555 3125 1645 3135
rect 1891 3125 2333 3135
rect 2595 3135 2605 3145
rect 2595 3125 2653 3135
rect 419 3105 797 3115
rect 1155 3105 1357 3115
rect 2355 3105 2813 3115
rect 3075 3105 3197 3115
rect 1155 3095 1165 3105
rect 1827 3095 2157 3105
rect 387 3085 461 3095
rect 1027 3085 1165 3095
rect 1331 3085 1837 3095
rect 2147 3085 2205 3095
rect 2355 3085 2413 3095
rect 2579 3085 2637 3095
rect 2707 3085 3149 3095
rect 803 3065 909 3075
rect 1379 3055 1389 3085
rect 2403 3075 2589 3085
rect 1587 3065 1661 3075
rect 1859 3065 1917 3075
rect 1987 3065 2237 3075
rect 1651 3055 1869 3065
rect 403 3045 621 3055
rect 1059 3045 1293 3055
rect 1347 3045 1389 3055
rect 2195 3045 2477 3055
rect 2659 3045 2877 3055
rect 1427 3035 1613 3045
rect 723 3025 813 3035
rect 1331 3025 1437 3035
rect 1603 3025 1837 3035
rect 1459 3005 1613 3015
rect 1731 3005 1885 3015
rect 1059 2985 1197 2995
rect 1219 2985 1437 2995
rect 1427 2975 1437 2985
rect 1587 2985 1725 2995
rect 2275 2985 2285 3045
rect 2675 3005 2925 3015
rect 2947 3005 3165 3015
rect 1587 2975 1597 2985
rect 1427 2965 1597 2975
rect 2083 2965 2317 2975
rect 2819 2965 2989 2975
rect 1763 2945 2045 2955
rect 2819 2945 2973 2955
rect 1763 2935 1773 2945
rect 1091 2925 1773 2935
rect 2035 2935 2045 2945
rect 2035 2925 2493 2935
rect 2627 2925 2797 2935
rect 2915 2925 2973 2935
rect 2787 2915 2925 2925
rect 1715 2905 1949 2915
rect 1491 2895 1677 2905
rect 1443 2885 1501 2895
rect 1667 2885 1757 2895
rect 1827 2885 2029 2895
rect 2531 2885 3021 2895
rect 915 2865 1245 2875
rect 1363 2865 1677 2875
rect 1731 2865 1869 2875
rect 2051 2865 2173 2875
rect 2371 2865 2525 2875
rect 1859 2855 2061 2865
rect 771 2825 973 2835
rect 1027 2815 1037 2855
rect 1523 2845 1821 2855
rect 1331 2835 1469 2845
rect 1171 2825 1341 2835
rect 1459 2825 1517 2835
rect 1555 2825 1789 2835
rect 1027 2805 1197 2815
rect 1363 2805 1661 2815
rect 643 2785 765 2795
rect 1219 2785 1805 2795
rect 1827 2785 1837 2835
rect 1859 2825 2029 2835
rect 2067 2825 2301 2835
rect 1859 2785 1869 2825
rect 2067 2815 2077 2825
rect 1891 2805 2077 2815
rect 2291 2815 2301 2825
rect 2339 2815 2349 2835
rect 2291 2805 2349 2815
rect 2371 2795 2381 2865
rect 2419 2845 2573 2855
rect 2643 2845 2797 2855
rect 2915 2845 3069 2855
rect 2467 2825 2541 2835
rect 2019 2785 2381 2795
rect 643 2775 653 2785
rect 2531 2775 2541 2825
rect 2563 2795 2573 2845
rect 2563 2785 2957 2795
rect 3091 2785 3325 2795
rect 595 2765 653 2775
rect 947 2765 1469 2775
rect 1923 2765 2109 2775
rect 2483 2765 2541 2775
rect 3027 2765 3165 2775
rect 1523 2755 1677 2765
rect 2163 2755 2445 2765
rect 547 2745 605 2755
rect 595 2735 605 2745
rect 787 2745 1069 2755
rect 1475 2745 1533 2755
rect 1667 2745 1933 2755
rect 2019 2745 2093 2755
rect 2115 2745 2173 2755
rect 2435 2745 2781 2755
rect 787 2735 797 2745
rect 1475 2735 1485 2745
rect 2115 2735 2125 2745
rect 595 2725 797 2735
rect 1219 2725 1485 2735
rect 1603 2725 1645 2735
rect 1811 2725 2125 2735
rect 2195 2725 2637 2735
rect 899 2705 1261 2715
rect 1395 2705 1629 2715
rect 1731 2705 1981 2715
rect 2035 2705 2749 2715
rect 2819 2705 3165 2715
rect 867 2685 1005 2695
rect 1027 2685 1181 2695
rect 1235 2685 1629 2695
rect 1779 2685 1965 2695
rect 1987 2685 2109 2695
rect 2211 2685 2509 2695
rect 2627 2685 2669 2695
rect 2211 2675 2221 2685
rect 579 2665 653 2675
rect 1379 2665 1453 2675
rect 1715 2665 1789 2675
rect 1859 2665 1917 2675
rect 2163 2665 2221 2675
rect 2259 2665 2317 2675
rect 979 2645 1197 2655
rect 1443 2645 1453 2665
rect 1907 2655 2173 2665
rect 2307 2655 2317 2665
rect 2659 2655 2669 2685
rect 2307 2645 2413 2655
rect 2467 2645 2637 2655
rect 2659 2645 2701 2655
rect 2835 2645 3165 2655
rect 979 2635 989 2645
rect 611 2625 989 2635
rect 1187 2635 1197 2645
rect 1619 2635 1773 2645
rect 1187 2625 1245 2635
rect 1363 2625 1629 2635
rect 1763 2625 1821 2635
rect 1859 2625 1917 2635
rect 1987 2625 2445 2635
rect 2483 2615 2749 2625
rect 2835 2615 2845 2645
rect 1011 2605 1101 2615
rect 1203 2605 1501 2615
rect 1651 2605 1965 2615
rect 2243 2605 2493 2615
rect 2739 2605 2845 2615
rect 3155 2615 3165 2645
rect 3155 2605 3357 2615
rect 691 2585 813 2595
rect 1347 2585 1437 2595
rect 1491 2585 1581 2595
rect 1827 2585 2013 2595
rect 2115 2585 2173 2595
rect 2435 2585 2701 2595
rect 803 2565 813 2585
rect 2163 2575 2445 2585
rect 2691 2575 2701 2585
rect 2867 2585 3133 2595
rect 2867 2575 2877 2585
rect 1747 2565 1933 2575
rect 2483 2565 2541 2575
rect 2691 2565 2877 2575
rect 1923 2555 2109 2565
rect 2483 2555 2493 2565
rect 1603 2545 1885 2555
rect 2099 2545 2493 2555
rect 1939 2525 2061 2535
rect 1107 2505 1565 2515
rect 1843 2505 1901 2515
rect 2083 2505 2781 2515
rect 1107 2495 1117 2505
rect 1059 2485 1117 2495
rect 1555 2495 1565 2505
rect 1891 2495 2093 2505
rect 1555 2485 1821 2495
rect 1811 2475 1821 2485
rect 2179 2485 2237 2495
rect 2179 2475 2189 2485
rect 739 2465 893 2475
rect 1811 2465 2189 2475
rect 739 2455 749 2465
rect 707 2445 749 2455
rect 883 2455 893 2465
rect 883 2445 1565 2455
rect 707 2425 717 2445
rect 2611 2425 2941 2435
rect 2611 2415 2621 2425
rect 723 2405 861 2415
rect 1539 2405 1933 2415
rect 2099 2405 2349 2415
rect 2387 2405 2621 2415
rect 2931 2415 2941 2425
rect 2931 2405 2989 2415
rect 2099 2395 2109 2405
rect 867 2385 1053 2395
rect 1203 2385 1309 2395
rect 1955 2385 2109 2395
rect 2339 2395 2349 2405
rect 2339 2385 2733 2395
rect 1843 2365 1981 2375
rect 2547 2365 3277 2375
rect 963 2345 1149 2355
rect 1187 2345 1357 2355
rect 2131 2345 2509 2355
rect 1187 2335 1197 2345
rect 899 2325 1197 2335
rect 1347 2335 1357 2345
rect 1347 2325 1405 2335
rect 1427 2325 1597 2335
rect 1987 2325 2253 2335
rect 611 2305 813 2315
rect 1027 2305 1533 2315
rect 2371 2305 2877 2315
rect 1107 2285 1229 2295
rect 1251 2285 1917 2295
rect 2211 2285 2301 2295
rect 2291 2275 2301 2285
rect 2419 2285 2477 2295
rect 2979 2285 3133 2295
rect 2419 2275 2429 2285
rect 1411 2265 1549 2275
rect 2291 2265 2429 2275
rect 819 2245 1261 2255
rect 1955 2245 2045 2255
rect 2083 2245 2253 2255
rect 1747 2225 1901 2235
rect 1011 2205 1181 2215
rect 1507 2205 1741 2215
rect 1843 2205 1901 2215
rect 2003 2205 2141 2215
rect 2339 2205 2445 2215
rect 1587 2185 1773 2195
rect 2227 2185 2333 2195
rect 2675 2185 3165 2195
rect 979 2165 1037 2175
rect 1027 2155 1037 2165
rect 1171 2165 1229 2175
rect 2355 2165 2589 2175
rect 1171 2155 1181 2165
rect 835 2145 973 2155
rect 1027 2145 1181 2155
rect 1315 2125 1405 2135
rect 1747 2105 2253 2115
rect 1747 2095 1757 2105
rect 1075 2085 1277 2095
rect 1075 2075 1085 2085
rect 1027 2065 1085 2075
rect 1267 2075 1277 2085
rect 1443 2085 1757 2095
rect 1443 2075 1453 2085
rect 1267 2065 1453 2075
rect 2243 2075 2253 2105
rect 2611 2085 2749 2095
rect 2243 2065 2525 2075
rect 739 2045 941 2055
rect 1283 2045 1341 2055
rect 1779 2045 1933 2055
rect 2099 2045 2221 2055
rect 2771 2045 2973 2055
rect 707 2025 813 2035
rect 899 2025 1261 2035
rect 1251 2015 1261 2025
rect 1379 2025 1677 2035
rect 1379 2015 1389 2025
rect 579 2005 861 2015
rect 1251 2005 1389 2015
rect 1475 2005 1581 2015
rect 2083 2005 2365 2015
rect 1539 1985 1645 1995
rect 1971 1985 2173 1995
rect 2755 1985 2909 1995
rect 899 1965 1021 1975
rect 1779 1965 1917 1975
rect 2147 1965 2493 1975
rect 2835 1965 3005 1975
rect 1203 1925 1341 1935
rect 1427 1925 2141 1935
rect 2403 1925 2653 1935
rect 1203 1915 1213 1925
rect 723 1905 861 1915
rect 723 1895 733 1905
rect 675 1885 733 1895
rect 851 1895 861 1905
rect 1091 1905 1213 1915
rect 1331 1915 1341 1925
rect 1331 1905 1981 1915
rect 1091 1895 1101 1905
rect 851 1885 1101 1895
rect 1235 1885 1613 1895
rect 1603 1875 1613 1885
rect 1763 1885 2077 1895
rect 2451 1885 2669 1895
rect 3235 1885 3405 1895
rect 1763 1875 1773 1885
rect 1603 1865 1773 1875
rect 1811 1865 1869 1875
rect 1859 1855 1869 1865
rect 2019 1865 2445 1875
rect 2019 1855 2029 1865
rect 595 1845 653 1855
rect 643 1835 653 1845
rect 771 1845 829 1855
rect 1123 1845 1245 1855
rect 1299 1845 1437 1855
rect 1859 1845 2029 1855
rect 2435 1855 2445 1865
rect 2435 1845 2621 1855
rect 771 1835 781 1845
rect 643 1825 781 1835
rect 1555 1825 1757 1835
rect 2067 1825 2125 1835
rect 2115 1815 2125 1825
rect 2275 1825 2477 1835
rect 2499 1825 2781 1835
rect 3171 1825 3437 1835
rect 2275 1815 2285 1825
rect 1603 1805 1773 1815
rect 2115 1805 2285 1815
rect 3363 1805 3485 1815
rect 1507 1785 1693 1795
rect 1827 1745 2141 1755
rect 1827 1735 1837 1745
rect 1219 1725 1373 1735
rect 1779 1725 1837 1735
rect 2131 1735 2141 1745
rect 2131 1725 2493 1735
rect 1411 1705 1565 1715
rect 1411 1695 1421 1705
rect 1235 1685 1421 1695
rect 1555 1695 1565 1705
rect 1555 1685 1773 1695
rect 1875 1685 1949 1695
rect 2019 1685 2109 1695
rect 3235 1685 3405 1695
rect 1139 1665 1229 1675
rect 1299 1665 1821 1675
rect 2147 1665 2349 1675
rect 1859 1655 2157 1665
rect 2339 1655 2349 1665
rect 1187 1645 1869 1655
rect 2339 1645 2477 1655
rect 2947 1645 3085 1655
rect 3363 1645 3485 1655
rect 563 1625 765 1635
rect 1267 1625 2093 1635
rect 2115 1625 2509 1635
rect 2083 1615 2093 1625
rect 1203 1605 1501 1615
rect 1523 1605 1597 1615
rect 2083 1605 2269 1615
rect 851 1585 989 1595
rect 1347 1575 1357 1605
rect 1443 1595 1453 1605
rect 1715 1595 1949 1605
rect 1443 1585 1725 1595
rect 1939 1585 2189 1595
rect 2339 1585 2349 1625
rect 2931 1605 3181 1615
rect 2499 1585 2637 1595
rect 3011 1585 3117 1595
rect 1299 1565 1357 1575
rect 1459 1565 1565 1575
rect 1747 1565 1869 1575
rect 2227 1565 2429 1575
rect 2467 1545 2525 1555
rect 2515 1535 2525 1545
rect 2643 1545 2781 1555
rect 3091 1545 3405 1555
rect 2643 1535 2653 1545
rect 595 1525 909 1535
rect 1315 1525 1821 1535
rect 2515 1525 2653 1535
rect 2771 1525 3069 1535
rect 1683 1505 1981 1515
rect 2099 1505 2397 1515
rect 2099 1495 2109 1505
rect 1235 1485 1661 1495
rect 1651 1475 1661 1485
rect 1875 1485 1933 1495
rect 2019 1485 2109 1495
rect 2387 1495 2397 1505
rect 2387 1485 2445 1495
rect 3027 1485 3293 1495
rect 1875 1475 1885 1485
rect 771 1465 1277 1475
rect 1651 1465 1885 1475
rect 1427 1445 1533 1455
rect 2131 1445 2589 1455
rect 739 1425 813 1435
rect 1779 1425 2109 1435
rect 2099 1415 2109 1425
rect 2515 1425 2573 1435
rect 851 1405 1005 1415
rect 1251 1405 1421 1415
rect 2099 1405 2253 1415
rect 851 1395 861 1405
rect 483 1385 861 1395
rect 995 1395 1005 1405
rect 2243 1395 2253 1405
rect 2515 1395 2525 1425
rect 995 1385 1053 1395
rect 2243 1385 2525 1395
rect 1155 1365 1805 1375
rect 1971 1365 2205 1375
rect 867 1345 1245 1355
rect 1075 1325 1133 1335
rect 1123 1315 1133 1325
rect 1331 1325 1389 1335
rect 2259 1325 2349 1335
rect 1331 1315 1341 1325
rect 1123 1305 1341 1315
rect 2243 1285 2429 1295
rect 2579 1285 2717 1295
rect 1731 1265 1853 1275
rect 1587 1245 1757 1255
rect 1987 1245 2109 1255
rect 2307 1245 2749 1255
rect 3443 1245 3565 1255
rect 963 1225 1021 1235
rect 1395 1225 1549 1235
rect 2355 1225 2557 1235
rect 2883 1225 3053 1235
rect 1395 1215 1405 1225
rect 1539 1215 1901 1225
rect 1075 1205 1405 1215
rect 1891 1205 1949 1215
rect 2115 1205 2301 1215
rect 2595 1205 2653 1215
rect 2643 1195 2653 1205
rect 2771 1205 2877 1215
rect 3411 1205 3581 1215
rect 2771 1195 2781 1205
rect 3411 1195 3421 1205
rect 755 1185 877 1195
rect 995 1185 1101 1195
rect 1571 1185 1965 1195
rect 2643 1185 2781 1195
rect 3123 1185 3261 1195
rect 3363 1185 3421 1195
rect 3571 1195 3581 1205
rect 3571 1185 3677 1195
rect 1427 1165 1629 1175
rect 2003 1165 2157 1175
rect 3379 1165 3453 1175
rect 1843 1155 2013 1165
rect 2147 1155 2157 1165
rect 3539 1155 3549 1175
rect 1683 1145 1853 1155
rect 2147 1145 2365 1155
rect 3539 1145 3565 1155
rect 835 1125 1165 1135
rect 1715 1125 2237 1135
rect 435 1105 573 1115
rect 1315 1105 1517 1115
rect 1667 1105 1789 1115
rect 2995 1105 3165 1115
rect 739 1085 1021 1095
rect 1123 1085 1229 1095
rect 1763 1085 2285 1095
rect 2611 1085 2733 1095
rect 2771 1085 2973 1095
rect 723 1045 829 1055
rect 1251 1035 1261 1075
rect 2195 1065 2525 1075
rect 1987 1045 2093 1055
rect 3555 1045 3565 1145
rect 499 1025 701 1035
rect 883 1025 941 1035
rect 1155 1025 1485 1035
rect 1699 1025 1789 1035
rect 2243 1025 2429 1035
rect 2579 1025 2669 1035
rect 3059 1025 3197 1035
rect 3283 1025 3389 1035
rect 691 1015 893 1025
rect 675 985 829 995
rect 819 975 829 985
rect 947 985 1005 995
rect 1299 985 1453 995
rect 1475 985 1965 995
rect 947 975 957 985
rect 819 965 957 975
rect 1635 945 1757 955
rect 451 925 781 935
rect 2147 925 2269 935
rect 3139 885 3293 895
rect 2515 865 3181 875
rect 595 845 765 855
rect 1459 845 2141 855
rect 3075 845 3213 855
rect 3267 845 3405 855
rect 947 825 1197 835
rect 2051 805 2509 815
rect 2819 805 2957 815
rect 467 785 813 795
rect 1171 785 1373 795
rect 1651 785 1853 795
rect 1891 785 2349 795
rect 2499 785 2509 805
rect 1651 775 1661 785
rect 723 765 1245 775
rect 1235 755 1245 765
rect 1395 765 1661 775
rect 1843 775 1853 785
rect 1843 765 2109 775
rect 1395 755 1405 765
rect 659 745 717 755
rect 899 745 1197 755
rect 1235 745 1405 755
rect 2339 755 2349 785
rect 2435 765 2605 775
rect 2339 745 2733 755
rect 707 735 909 745
rect 1619 725 1965 735
rect 2675 725 2909 735
rect 787 705 1181 715
rect 1379 705 1645 715
rect 2227 705 2397 715
rect 2419 705 2701 715
rect 2691 695 2701 705
rect 627 685 765 695
rect 1411 685 1469 695
rect 1459 675 1469 685
rect 1619 685 1901 695
rect 1939 685 2525 695
rect 2691 685 2845 695
rect 3523 685 3581 695
rect 1619 675 1629 685
rect 1459 665 1629 675
rect 1891 675 1901 685
rect 1891 665 2125 675
rect 2387 665 2445 675
rect 3299 665 3357 675
rect 2115 655 2397 665
rect 547 645 685 655
rect 723 645 973 655
rect 1379 625 1613 635
rect 1891 625 1949 635
rect 1939 615 1949 625
rect 2115 625 2173 635
rect 2275 625 2333 635
rect 2115 615 2125 625
rect 1939 605 2125 615
rect 2323 615 2333 625
rect 2451 625 2749 635
rect 3299 625 3309 665
rect 3331 625 3597 635
rect 2451 615 2461 625
rect 2323 605 2461 615
rect 2499 605 2621 615
rect 339 585 685 595
rect 2611 585 2765 595
rect 723 565 941 575
rect 2563 565 2637 575
rect 3251 485 3581 495
rect 1507 465 1677 475
rect 1507 435 1517 465
rect 1667 455 1677 465
rect 1667 445 1725 455
rect 1955 445 2045 455
rect 2339 445 2541 455
rect 3267 445 3517 455
rect 675 425 1517 435
rect 3091 425 3245 435
rect 3443 425 3501 435
rect 3235 415 3453 425
rect 1523 405 1837 415
rect 1923 405 2029 415
rect 2179 385 2349 395
rect 2899 385 3021 395
rect 3171 385 3229 395
rect 3443 385 3629 395
rect 3171 375 3181 385
rect 1667 365 1869 375
rect 2947 365 3181 375
rect 3219 365 3325 375
rect 2531 345 2925 355
rect 2835 325 3165 335
rect 1331 285 1517 295
rect 2723 285 3069 295
rect 1475 265 1757 275
rect 1315 225 1597 235
rect 2643 225 3085 235
rect 2627 185 2845 195
use AND2X2  AND2X2_0
timestamp 1090541974
transform 1 0 2816 0 -1 1940
box -16 -6 80 210
use AND2X2  AND2X2_1
timestamp 1090541974
transform 1 0 592 0 1 1140
box -16 -6 80 210
use AND2X2  AND2X2_2
timestamp 1090541974
transform 1 0 1056 0 -1 1140
box -16 -6 80 210
use AND2X2  AND2X2_3
timestamp 1090541974
transform 1 0 1232 0 1 1140
box -16 -6 80 210
use AOI21X1  AOI21X1_0
timestamp 1090541997
transform 1 0 704 0 1 740
box -14 -6 78 210
use AOI21X1  AOI21X1_1
timestamp 1090541997
transform 1 0 736 0 -1 1540
box -14 -6 78 210
use AOI21X1  AOI21X1_2
timestamp 1090541997
transform 1 0 928 0 1 740
box -14 -6 78 210
use AOI21X1  AOI21X1_3
timestamp 1090541997
transform 1 0 1440 0 1 340
box -14 -6 78 210
use AOI21X1  AOI21X1_4
timestamp 1090541997
transform 1 0 1680 0 -1 340
box -14 -6 78 210
use AOI22X1  AOI22X1_0
timestamp 1053022145
transform 1 0 2432 0 1 740
box -16 -6 92 210
use AOI22X1  AOI22X1_1
timestamp 1053022145
transform 1 0 2080 0 -1 740
box -16 -6 92 210
use AOI22X1  AOI22X1_2
timestamp 1053022145
transform 1 0 1888 0 -1 740
box -16 -6 92 210
use AOI22X1  AOI22X1_3
timestamp 1053022145
transform 1 0 2576 0 -1 1140
box -16 -6 92 210
use AOI22X1  AOI22X1_4
timestamp 1053022145
transform 1 0 1840 0 1 3140
box -16 -6 92 210
use AOI22X1  AOI22X1_5
timestamp 1053022145
transform 1 0 1728 0 -1 2740
box -16 -6 92 210
use AOI22X1  AOI22X1_6
timestamp 1053022145
transform 1 0 1824 0 -1 2740
box -16 -6 92 210
use AOI22X1  AOI22X1_7
timestamp 1053022145
transform 1 0 1968 0 1 2340
box -16 -6 92 210
use AOI22X1  AOI22X1_8
timestamp 1053022145
transform 1 0 1824 0 1 2340
box -16 -6 92 210
use DFFNEGX1  DFFNEGX1_0
timestamp 1052851797
transform 1 0 2752 0 -1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_1
timestamp 1052851797
transform 1 0 2704 0 1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_2
timestamp 1052851797
transform 1 0 2944 0 -1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_3
timestamp 1052851797
transform 1 0 2960 0 1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_4
timestamp 1052851797
transform 1 0 2944 0 -1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_5
timestamp 1052851797
transform 1 0 3040 0 -1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_6
timestamp 1052851797
transform 1 0 2832 0 1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_7
timestamp 1052851797
transform 1 0 2992 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_8
timestamp 1052851797
transform 1 0 2528 0 1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_9
timestamp 1052851797
transform 1 0 1840 0 1 340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_10
timestamp 1052851797
transform 1 0 1872 0 1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_11
timestamp 1052851797
transform 1 0 2160 0 1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_12
timestamp 1052851797
transform 1 0 2336 0 1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_13
timestamp 1052851797
transform 1 0 1152 0 1 340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_14
timestamp 1052851797
transform 1 0 320 0 -1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_15
timestamp 1052851797
transform 1 0 656 0 1 340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_16
timestamp 1052851797
transform 1 0 320 0 -1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_17
timestamp 1052851797
transform 1 0 2560 0 1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_18
timestamp 1052851797
transform 1 0 2592 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_19
timestamp 1052851797
transform 1 0 1792 0 1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_20
timestamp 1052851797
transform 1 0 1440 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_21
timestamp 1052851797
transform 1 0 1776 0 1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_22
timestamp 1052851797
transform 1 0 1664 0 1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_23
timestamp 1052851797
transform 1 0 2336 0 -1 1140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_24
timestamp 1052851797
transform 1 0 2240 0 -1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_25
timestamp 1052851797
transform 1 0 1280 0 1 1540
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_26
timestamp 1052851797
transform 1 0 1040 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_27
timestamp 1052851797
transform 1 0 1952 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_28
timestamp 1052851797
transform 1 0 656 0 -1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_29
timestamp 1052851797
transform 1 0 1936 0 -1 2340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_30
timestamp 1052851797
transform 1 0 1136 0 1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_31
timestamp 1052851797
transform 1 0 1360 0 1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_32
timestamp 1052851797
transform 1 0 2144 0 1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_33
timestamp 1052851797
transform 1 0 2912 0 -1 2740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_34
timestamp 1052851797
transform 1 0 672 0 -1 2740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_35
timestamp 1052851797
transform 1 0 784 0 1 2340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_36
timestamp 1052851797
transform 1 0 3136 0 -1 2740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_37
timestamp 1052851797
transform 1 0 2032 0 1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_38
timestamp 1052851797
transform 1 0 2752 0 1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_39
timestamp 1052851797
transform 1 0 2976 0 1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_40
timestamp 1052851797
transform 1 0 2416 0 1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_41
timestamp 1052851797
transform 1 0 2960 0 -1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_42
timestamp 1052851797
transform 1 0 832 0 -1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_43
timestamp 1052851797
transform 1 0 1056 0 1 3140
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_44
timestamp 1052851797
transform 1 0 2800 0 1 2740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_45
timestamp 1052851797
transform 1 0 2656 0 1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_46
timestamp 1052851797
transform 1 0 592 0 -1 2340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_47
timestamp 1052851797
transform 1 0 944 0 1 1940
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_48
timestamp 1052851797
transform 1 0 3056 0 -1 2340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_49
timestamp 1052851797
transform 1 0 1648 0 1 340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_50
timestamp 1052851797
transform 1 0 1136 0 -1 340
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_51
timestamp 1052851797
transform 1 0 1424 0 -1 740
box -16 -6 208 210
use DFFNEGX1  DFFNEGX1_52
timestamp 1052851797
transform 1 0 1616 0 -1 740
box -16 -6 208 210
use FILL  FILL_0
timestamp 1018054153
transform 1 0 3664 0 -1 3540
box -16 -6 32 210
use FILL  FILL_1
timestamp 1018054153
transform 1 0 3648 0 -1 3540
box -16 -6 32 210
use FILL  FILL_2
timestamp 1018054153
transform 1 0 3632 0 -1 3540
box -16 -6 32 210
use FILL  FILL_3
timestamp 1018054153
transform 1 0 3616 0 -1 3540
box -16 -6 32 210
use FILL  FILL_4
timestamp 1018054153
transform 1 0 3600 0 -1 3540
box -16 -6 32 210
use FILL  FILL_5
timestamp 1018054153
transform 1 0 3584 0 -1 3540
box -16 -6 32 210
use FILL  FILL_6
timestamp 1018054153
transform 1 0 3568 0 -1 3540
box -16 -6 32 210
use FILL  FILL_7
timestamp 1018054153
transform 1 0 3552 0 -1 3540
box -16 -6 32 210
use FILL  FILL_8
timestamp 1018054153
transform 1 0 3536 0 -1 3540
box -16 -6 32 210
use FILL  FILL_9
timestamp 1018054153
transform 1 0 3520 0 -1 3540
box -16 -6 32 210
use FILL  FILL_10
timestamp 1018054153
transform 1 0 3504 0 -1 3540
box -16 -6 32 210
use FILL  FILL_11
timestamp 1018054153
transform 1 0 3488 0 -1 3540
box -16 -6 32 210
use FILL  FILL_12
timestamp 1018054153
transform 1 0 3472 0 -1 3540
box -16 -6 32 210
use FILL  FILL_13
timestamp 1018054153
transform 1 0 3456 0 -1 3540
box -16 -6 32 210
use FILL  FILL_14
timestamp 1018054153
transform 1 0 3440 0 -1 3540
box -16 -6 32 210
use FILL  FILL_15
timestamp 1018054153
transform 1 0 3424 0 -1 3540
box -16 -6 32 210
use FILL  FILL_16
timestamp 1018054153
transform 1 0 3408 0 -1 3540
box -16 -6 32 210
use FILL  FILL_17
timestamp 1018054153
transform 1 0 3392 0 -1 3540
box -16 -6 32 210
use FILL  FILL_18
timestamp 1018054153
transform 1 0 3376 0 -1 3540
box -16 -6 32 210
use FILL  FILL_19
timestamp 1018054153
transform 1 0 3360 0 -1 3540
box -16 -6 32 210
use FILL  FILL_20
timestamp 1018054153
transform 1 0 3344 0 -1 3540
box -16 -6 32 210
use FILL  FILL_21
timestamp 1018054153
transform 1 0 3328 0 -1 3540
box -16 -6 32 210
use FILL  FILL_22
timestamp 1018054153
transform 1 0 3312 0 -1 3540
box -16 -6 32 210
use FILL  FILL_23
timestamp 1018054153
transform 1 0 3296 0 -1 3540
box -16 -6 32 210
use FILL  FILL_24
timestamp 1018054153
transform 1 0 3280 0 -1 3540
box -16 -6 32 210
use FILL  FILL_25
timestamp 1018054153
transform 1 0 3264 0 -1 3540
box -16 -6 32 210
use FILL  FILL_26
timestamp 1018054153
transform 1 0 3248 0 -1 3540
box -16 -6 32 210
use FILL  FILL_27
timestamp 1018054153
transform 1 0 3200 0 -1 3540
box -16 -6 32 210
use FILL  FILL_28
timestamp 1018054153
transform 1 0 3184 0 -1 3540
box -16 -6 32 210
use FILL  FILL_29
timestamp 1018054153
transform 1 0 3168 0 -1 3540
box -16 -6 32 210
use FILL  FILL_30
timestamp 1018054153
transform 1 0 3152 0 -1 3540
box -16 -6 32 210
use FILL  FILL_31
timestamp 1018054153
transform 1 0 3024 0 -1 3540
box -16 -6 32 210
use FILL  FILL_32
timestamp 1018054153
transform 1 0 3008 0 -1 3540
box -16 -6 32 210
use FILL  FILL_33
timestamp 1018054153
transform 1 0 2992 0 -1 3540
box -16 -6 32 210
use FILL  FILL_34
timestamp 1018054153
transform 1 0 2976 0 -1 3540
box -16 -6 32 210
use FILL  FILL_35
timestamp 1018054153
transform 1 0 2960 0 -1 3540
box -16 -6 32 210
use FILL  FILL_36
timestamp 1018054153
transform 1 0 2944 0 -1 3540
box -16 -6 32 210
use FILL  FILL_37
timestamp 1018054153
transform 1 0 2928 0 -1 3540
box -16 -6 32 210
use FILL  FILL_38
timestamp 1018054153
transform 1 0 2912 0 -1 3540
box -16 -6 32 210
use FILL  FILL_39
timestamp 1018054153
transform 1 0 2896 0 -1 3540
box -16 -6 32 210
use FILL  FILL_40
timestamp 1018054153
transform 1 0 2768 0 -1 3540
box -16 -6 32 210
use FILL  FILL_41
timestamp 1018054153
transform 1 0 2752 0 -1 3540
box -16 -6 32 210
use FILL  FILL_42
timestamp 1018054153
transform 1 0 2736 0 -1 3540
box -16 -6 32 210
use FILL  FILL_43
timestamp 1018054153
transform 1 0 2688 0 -1 3540
box -16 -6 32 210
use FILL  FILL_44
timestamp 1018054153
transform 1 0 2672 0 -1 3540
box -16 -6 32 210
use FILL  FILL_45
timestamp 1018054153
transform 1 0 2656 0 -1 3540
box -16 -6 32 210
use FILL  FILL_46
timestamp 1018054153
transform 1 0 2640 0 -1 3540
box -16 -6 32 210
use FILL  FILL_47
timestamp 1018054153
transform 1 0 2624 0 -1 3540
box -16 -6 32 210
use FILL  FILL_48
timestamp 1018054153
transform 1 0 2608 0 -1 3540
box -16 -6 32 210
use FILL  FILL_49
timestamp 1018054153
transform 1 0 2592 0 -1 3540
box -16 -6 32 210
use FILL  FILL_50
timestamp 1018054153
transform 1 0 2576 0 -1 3540
box -16 -6 32 210
use FILL  FILL_51
timestamp 1018054153
transform 1 0 2560 0 -1 3540
box -16 -6 32 210
use FILL  FILL_52
timestamp 1018054153
transform 1 0 2432 0 -1 3540
box -16 -6 32 210
use FILL  FILL_53
timestamp 1018054153
transform 1 0 2416 0 -1 3540
box -16 -6 32 210
use FILL  FILL_54
timestamp 1018054153
transform 1 0 2400 0 -1 3540
box -16 -6 32 210
use FILL  FILL_55
timestamp 1018054153
transform 1 0 2384 0 -1 3540
box -16 -6 32 210
use FILL  FILL_56
timestamp 1018054153
transform 1 0 2368 0 -1 3540
box -16 -6 32 210
use FILL  FILL_57
timestamp 1018054153
transform 1 0 2352 0 -1 3540
box -16 -6 32 210
use FILL  FILL_58
timestamp 1018054153
transform 1 0 2336 0 -1 3540
box -16 -6 32 210
use FILL  FILL_59
timestamp 1018054153
transform 1 0 2320 0 -1 3540
box -16 -6 32 210
use FILL  FILL_60
timestamp 1018054153
transform 1 0 2304 0 -1 3540
box -16 -6 32 210
use FILL  FILL_61
timestamp 1018054153
transform 1 0 2288 0 -1 3540
box -16 -6 32 210
use FILL  FILL_62
timestamp 1018054153
transform 1 0 2272 0 -1 3540
box -16 -6 32 210
use FILL  FILL_63
timestamp 1018054153
transform 1 0 2256 0 -1 3540
box -16 -6 32 210
use FILL  FILL_64
timestamp 1018054153
transform 1 0 2240 0 -1 3540
box -16 -6 32 210
use FILL  FILL_65
timestamp 1018054153
transform 1 0 2224 0 -1 3540
box -16 -6 32 210
use FILL  FILL_66
timestamp 1018054153
transform 1 0 2096 0 -1 3540
box -16 -6 32 210
use FILL  FILL_67
timestamp 1018054153
transform 1 0 2080 0 -1 3540
box -16 -6 32 210
use FILL  FILL_68
timestamp 1018054153
transform 1 0 2064 0 -1 3540
box -16 -6 32 210
use FILL  FILL_69
timestamp 1018054153
transform 1 0 2048 0 -1 3540
box -16 -6 32 210
use FILL  FILL_70
timestamp 1018054153
transform 1 0 2032 0 -1 3540
box -16 -6 32 210
use FILL  FILL_71
timestamp 1018054153
transform 1 0 2016 0 -1 3540
box -16 -6 32 210
use FILL  FILL_72
timestamp 1018054153
transform 1 0 2000 0 -1 3540
box -16 -6 32 210
use FILL  FILL_73
timestamp 1018054153
transform 1 0 1984 0 -1 3540
box -16 -6 32 210
use FILL  FILL_74
timestamp 1018054153
transform 1 0 1968 0 -1 3540
box -16 -6 32 210
use FILL  FILL_75
timestamp 1018054153
transform 1 0 1952 0 -1 3540
box -16 -6 32 210
use FILL  FILL_76
timestamp 1018054153
transform 1 0 1824 0 -1 3540
box -16 -6 32 210
use FILL  FILL_77
timestamp 1018054153
transform 1 0 1808 0 -1 3540
box -16 -6 32 210
use FILL  FILL_78
timestamp 1018054153
transform 1 0 1568 0 -1 3540
box -16 -6 32 210
use FILL  FILL_79
timestamp 1018054153
transform 1 0 1552 0 -1 3540
box -16 -6 32 210
use FILL  FILL_80
timestamp 1018054153
transform 1 0 1536 0 -1 3540
box -16 -6 32 210
use FILL  FILL_81
timestamp 1018054153
transform 1 0 1520 0 -1 3540
box -16 -6 32 210
use FILL  FILL_82
timestamp 1018054153
transform 1 0 1504 0 -1 3540
box -16 -6 32 210
use FILL  FILL_83
timestamp 1018054153
transform 1 0 1456 0 -1 3540
box -16 -6 32 210
use FILL  FILL_84
timestamp 1018054153
transform 1 0 1440 0 -1 3540
box -16 -6 32 210
use FILL  FILL_85
timestamp 1018054153
transform 1 0 1424 0 -1 3540
box -16 -6 32 210
use FILL  FILL_86
timestamp 1018054153
transform 1 0 1408 0 -1 3540
box -16 -6 32 210
use FILL  FILL_87
timestamp 1018054153
transform 1 0 1392 0 -1 3540
box -16 -6 32 210
use FILL  FILL_88
timestamp 1018054153
transform 1 0 1376 0 -1 3540
box -16 -6 32 210
use FILL  FILL_89
timestamp 1018054153
transform 1 0 1360 0 -1 3540
box -16 -6 32 210
use FILL  FILL_90
timestamp 1018054153
transform 1 0 1344 0 -1 3540
box -16 -6 32 210
use FILL  FILL_91
timestamp 1018054153
transform 1 0 1328 0 -1 3540
box -16 -6 32 210
use FILL  FILL_92
timestamp 1018054153
transform 1 0 1312 0 -1 3540
box -16 -6 32 210
use FILL  FILL_93
timestamp 1018054153
transform 1 0 1296 0 -1 3540
box -16 -6 32 210
use FILL  FILL_94
timestamp 1018054153
transform 1 0 1280 0 -1 3540
box -16 -6 32 210
use FILL  FILL_95
timestamp 1018054153
transform 1 0 1264 0 -1 3540
box -16 -6 32 210
use FILL  FILL_96
timestamp 1018054153
transform 1 0 1248 0 -1 3540
box -16 -6 32 210
use FILL  FILL_97
timestamp 1018054153
transform 1 0 1120 0 -1 3540
box -16 -6 32 210
use FILL  FILL_98
timestamp 1018054153
transform 1 0 1104 0 -1 3540
box -16 -6 32 210
use FILL  FILL_99
timestamp 1018054153
transform 1 0 1088 0 -1 3540
box -16 -6 32 210
use FILL  FILL_100
timestamp 1018054153
transform 1 0 1072 0 -1 3540
box -16 -6 32 210
use FILL  FILL_101
timestamp 1018054153
transform 1 0 1056 0 -1 3540
box -16 -6 32 210
use FILL  FILL_102
timestamp 1018054153
transform 1 0 1040 0 -1 3540
box -16 -6 32 210
use FILL  FILL_103
timestamp 1018054153
transform 1 0 1024 0 -1 3540
box -16 -6 32 210
use FILL  FILL_104
timestamp 1018054153
transform 1 0 1008 0 -1 3540
box -16 -6 32 210
use FILL  FILL_105
timestamp 1018054153
transform 1 0 992 0 -1 3540
box -16 -6 32 210
use FILL  FILL_106
timestamp 1018054153
transform 1 0 976 0 -1 3540
box -16 -6 32 210
use FILL  FILL_107
timestamp 1018054153
transform 1 0 960 0 -1 3540
box -16 -6 32 210
use FILL  FILL_108
timestamp 1018054153
transform 1 0 944 0 -1 3540
box -16 -6 32 210
use FILL  FILL_109
timestamp 1018054153
transform 1 0 928 0 -1 3540
box -16 -6 32 210
use FILL  FILL_110
timestamp 1018054153
transform 1 0 912 0 -1 3540
box -16 -6 32 210
use FILL  FILL_111
timestamp 1018054153
transform 1 0 896 0 -1 3540
box -16 -6 32 210
use FILL  FILL_112
timestamp 1018054153
transform 1 0 880 0 -1 3540
box -16 -6 32 210
use FILL  FILL_113
timestamp 1018054153
transform 1 0 864 0 -1 3540
box -16 -6 32 210
use FILL  FILL_114
timestamp 1018054153
transform 1 0 848 0 -1 3540
box -16 -6 32 210
use FILL  FILL_115
timestamp 1018054153
transform 1 0 832 0 -1 3540
box -16 -6 32 210
use FILL  FILL_116
timestamp 1018054153
transform 1 0 816 0 -1 3540
box -16 -6 32 210
use FILL  FILL_117
timestamp 1018054153
transform 1 0 800 0 -1 3540
box -16 -6 32 210
use FILL  FILL_118
timestamp 1018054153
transform 1 0 784 0 -1 3540
box -16 -6 32 210
use FILL  FILL_119
timestamp 1018054153
transform 1 0 768 0 -1 3540
box -16 -6 32 210
use FILL  FILL_120
timestamp 1018054153
transform 1 0 752 0 -1 3540
box -16 -6 32 210
use FILL  FILL_121
timestamp 1018054153
transform 1 0 736 0 -1 3540
box -16 -6 32 210
use FILL  FILL_122
timestamp 1018054153
transform 1 0 720 0 -1 3540
box -16 -6 32 210
use FILL  FILL_123
timestamp 1018054153
transform 1 0 704 0 -1 3540
box -16 -6 32 210
use FILL  FILL_124
timestamp 1018054153
transform 1 0 688 0 -1 3540
box -16 -6 32 210
use FILL  FILL_125
timestamp 1018054153
transform 1 0 672 0 -1 3540
box -16 -6 32 210
use FILL  FILL_126
timestamp 1018054153
transform 1 0 656 0 -1 3540
box -16 -6 32 210
use FILL  FILL_127
timestamp 1018054153
transform 1 0 640 0 -1 3540
box -16 -6 32 210
use FILL  FILL_128
timestamp 1018054153
transform 1 0 624 0 -1 3540
box -16 -6 32 210
use FILL  FILL_129
timestamp 1018054153
transform 1 0 608 0 -1 3540
box -16 -6 32 210
use FILL  FILL_130
timestamp 1018054153
transform 1 0 592 0 -1 3540
box -16 -6 32 210
use FILL  FILL_131
timestamp 1018054153
transform 1 0 576 0 -1 3540
box -16 -6 32 210
use FILL  FILL_132
timestamp 1018054153
transform 1 0 560 0 -1 3540
box -16 -6 32 210
use FILL  FILL_133
timestamp 1018054153
transform 1 0 544 0 -1 3540
box -16 -6 32 210
use FILL  FILL_134
timestamp 1018054153
transform 1 0 528 0 -1 3540
box -16 -6 32 210
use FILL  FILL_135
timestamp 1018054153
transform 1 0 512 0 -1 3540
box -16 -6 32 210
use FILL  FILL_136
timestamp 1018054153
transform 1 0 496 0 -1 3540
box -16 -6 32 210
use FILL  FILL_137
timestamp 1018054153
transform 1 0 480 0 -1 3540
box -16 -6 32 210
use FILL  FILL_138
timestamp 1018054153
transform 1 0 464 0 -1 3540
box -16 -6 32 210
use FILL  FILL_139
timestamp 1018054153
transform 1 0 448 0 -1 3540
box -16 -6 32 210
use FILL  FILL_140
timestamp 1018054153
transform 1 0 432 0 -1 3540
box -16 -6 32 210
use FILL  FILL_141
timestamp 1018054153
transform 1 0 416 0 -1 3540
box -16 -6 32 210
use FILL  FILL_142
timestamp 1018054153
transform 1 0 400 0 -1 3540
box -16 -6 32 210
use FILL  FILL_143
timestamp 1018054153
transform 1 0 384 0 -1 3540
box -16 -6 32 210
use FILL  FILL_144
timestamp 1018054153
transform 1 0 368 0 -1 3540
box -16 -6 32 210
use FILL  FILL_145
timestamp 1018054153
transform 1 0 352 0 -1 3540
box -16 -6 32 210
use FILL  FILL_146
timestamp 1018054153
transform 1 0 336 0 -1 3540
box -16 -6 32 210
use FILL  FILL_147
timestamp 1018054153
transform 1 0 320 0 -1 3540
box -16 -6 32 210
use FILL  FILL_148
timestamp 1018054153
transform 1 0 304 0 -1 3540
box -16 -6 32 210
use FILL  FILL_149
timestamp 1018054153
transform 1 0 288 0 -1 3540
box -16 -6 32 210
use FILL  FILL_150
timestamp 1018054153
transform 1 0 272 0 -1 3540
box -16 -6 32 210
use FILL  FILL_151
timestamp 1018054153
transform 1 0 256 0 -1 3540
box -16 -6 32 210
use FILL  FILL_152
timestamp 1018054153
transform 1 0 240 0 -1 3540
box -16 -6 32 210
use FILL  FILL_153
timestamp 1018054153
transform 1 0 224 0 -1 3540
box -16 -6 32 210
use FILL  FILL_154
timestamp 1018054153
transform 1 0 208 0 -1 3540
box -16 -6 32 210
use FILL  FILL_155
timestamp 1018054153
transform 1 0 192 0 -1 3540
box -16 -6 32 210
use FILL  FILL_156
timestamp 1018054153
transform 1 0 176 0 -1 3540
box -16 -6 32 210
use FILL  FILL_157
timestamp 1018054153
transform 1 0 160 0 -1 3540
box -16 -6 32 210
use FILL  FILL_158
timestamp 1018054153
transform 1 0 144 0 -1 3540
box -16 -6 32 210
use FILL  FILL_159
timestamp 1018054153
transform 1 0 3664 0 1 3140
box -16 -6 32 210
use FILL  FILL_160
timestamp 1018054153
transform 1 0 3648 0 1 3140
box -16 -6 32 210
use FILL  FILL_161
timestamp 1018054153
transform 1 0 3632 0 1 3140
box -16 -6 32 210
use FILL  FILL_162
timestamp 1018054153
transform 1 0 3616 0 1 3140
box -16 -6 32 210
use FILL  FILL_163
timestamp 1018054153
transform 1 0 3600 0 1 3140
box -16 -6 32 210
use FILL  FILL_164
timestamp 1018054153
transform 1 0 3584 0 1 3140
box -16 -6 32 210
use FILL  FILL_165
timestamp 1018054153
transform 1 0 3568 0 1 3140
box -16 -6 32 210
use FILL  FILL_166
timestamp 1018054153
transform 1 0 3552 0 1 3140
box -16 -6 32 210
use FILL  FILL_167
timestamp 1018054153
transform 1 0 3536 0 1 3140
box -16 -6 32 210
use FILL  FILL_168
timestamp 1018054153
transform 1 0 3520 0 1 3140
box -16 -6 32 210
use FILL  FILL_169
timestamp 1018054153
transform 1 0 3504 0 1 3140
box -16 -6 32 210
use FILL  FILL_170
timestamp 1018054153
transform 1 0 3488 0 1 3140
box -16 -6 32 210
use FILL  FILL_171
timestamp 1018054153
transform 1 0 3472 0 1 3140
box -16 -6 32 210
use FILL  FILL_172
timestamp 1018054153
transform 1 0 3456 0 1 3140
box -16 -6 32 210
use FILL  FILL_173
timestamp 1018054153
transform 1 0 3440 0 1 3140
box -16 -6 32 210
use FILL  FILL_174
timestamp 1018054153
transform 1 0 3424 0 1 3140
box -16 -6 32 210
use FILL  FILL_175
timestamp 1018054153
transform 1 0 3408 0 1 3140
box -16 -6 32 210
use FILL  FILL_176
timestamp 1018054153
transform 1 0 3392 0 1 3140
box -16 -6 32 210
use FILL  FILL_177
timestamp 1018054153
transform 1 0 3376 0 1 3140
box -16 -6 32 210
use FILL  FILL_178
timestamp 1018054153
transform 1 0 3360 0 1 3140
box -16 -6 32 210
use FILL  FILL_179
timestamp 1018054153
transform 1 0 3344 0 1 3140
box -16 -6 32 210
use FILL  FILL_180
timestamp 1018054153
transform 1 0 3328 0 1 3140
box -16 -6 32 210
use FILL  FILL_181
timestamp 1018054153
transform 1 0 3312 0 1 3140
box -16 -6 32 210
use FILL  FILL_182
timestamp 1018054153
transform 1 0 3296 0 1 3140
box -16 -6 32 210
use FILL  FILL_183
timestamp 1018054153
transform 1 0 3280 0 1 3140
box -16 -6 32 210
use FILL  FILL_184
timestamp 1018054153
transform 1 0 3264 0 1 3140
box -16 -6 32 210
use FILL  FILL_185
timestamp 1018054153
transform 1 0 3248 0 1 3140
box -16 -6 32 210
use FILL  FILL_186
timestamp 1018054153
transform 1 0 3232 0 1 3140
box -16 -6 32 210
use FILL  FILL_187
timestamp 1018054153
transform 1 0 3216 0 1 3140
box -16 -6 32 210
use FILL  FILL_188
timestamp 1018054153
transform 1 0 3200 0 1 3140
box -16 -6 32 210
use FILL  FILL_189
timestamp 1018054153
transform 1 0 3184 0 1 3140
box -16 -6 32 210
use FILL  FILL_190
timestamp 1018054153
transform 1 0 3168 0 1 3140
box -16 -6 32 210
use FILL  FILL_191
timestamp 1018054153
transform 1 0 2960 0 1 3140
box -16 -6 32 210
use FILL  FILL_192
timestamp 1018054153
transform 1 0 2944 0 1 3140
box -16 -6 32 210
use FILL  FILL_193
timestamp 1018054153
transform 1 0 1680 0 1 3140
box -16 -6 32 210
use FILL  FILL_194
timestamp 1018054153
transform 1 0 1664 0 1 3140
box -16 -6 32 210
use FILL  FILL_195
timestamp 1018054153
transform 1 0 1648 0 1 3140
box -16 -6 32 210
use FILL  FILL_196
timestamp 1018054153
transform 1 0 1344 0 1 3140
box -16 -6 32 210
use FILL  FILL_197
timestamp 1018054153
transform 1 0 1328 0 1 3140
box -16 -6 32 210
use FILL  FILL_198
timestamp 1018054153
transform 1 0 1312 0 1 3140
box -16 -6 32 210
use FILL  FILL_199
timestamp 1018054153
transform 1 0 1296 0 1 3140
box -16 -6 32 210
use FILL  FILL_200
timestamp 1018054153
transform 1 0 1280 0 1 3140
box -16 -6 32 210
use FILL  FILL_201
timestamp 1018054153
transform 1 0 1040 0 1 3140
box -16 -6 32 210
use FILL  FILL_202
timestamp 1018054153
transform 1 0 848 0 1 3140
box -16 -6 32 210
use FILL  FILL_203
timestamp 1018054153
transform 1 0 832 0 1 3140
box -16 -6 32 210
use FILL  FILL_204
timestamp 1018054153
transform 1 0 736 0 1 3140
box -16 -6 32 210
use FILL  FILL_205
timestamp 1018054153
transform 1 0 720 0 1 3140
box -16 -6 32 210
use FILL  FILL_206
timestamp 1018054153
transform 1 0 704 0 1 3140
box -16 -6 32 210
use FILL  FILL_207
timestamp 1018054153
transform 1 0 688 0 1 3140
box -16 -6 32 210
use FILL  FILL_208
timestamp 1018054153
transform 1 0 528 0 1 3140
box -16 -6 32 210
use FILL  FILL_209
timestamp 1018054153
transform 1 0 512 0 1 3140
box -16 -6 32 210
use FILL  FILL_210
timestamp 1018054153
transform 1 0 496 0 1 3140
box -16 -6 32 210
use FILL  FILL_211
timestamp 1018054153
transform 1 0 480 0 1 3140
box -16 -6 32 210
use FILL  FILL_212
timestamp 1018054153
transform 1 0 464 0 1 3140
box -16 -6 32 210
use FILL  FILL_213
timestamp 1018054153
transform 1 0 448 0 1 3140
box -16 -6 32 210
use FILL  FILL_214
timestamp 1018054153
transform 1 0 432 0 1 3140
box -16 -6 32 210
use FILL  FILL_215
timestamp 1018054153
transform 1 0 416 0 1 3140
box -16 -6 32 210
use FILL  FILL_216
timestamp 1018054153
transform 1 0 400 0 1 3140
box -16 -6 32 210
use FILL  FILL_217
timestamp 1018054153
transform 1 0 384 0 1 3140
box -16 -6 32 210
use FILL  FILL_218
timestamp 1018054153
transform 1 0 368 0 1 3140
box -16 -6 32 210
use FILL  FILL_219
timestamp 1018054153
transform 1 0 352 0 1 3140
box -16 -6 32 210
use FILL  FILL_220
timestamp 1018054153
transform 1 0 336 0 1 3140
box -16 -6 32 210
use FILL  FILL_221
timestamp 1018054153
transform 1 0 320 0 1 3140
box -16 -6 32 210
use FILL  FILL_222
timestamp 1018054153
transform 1 0 304 0 1 3140
box -16 -6 32 210
use FILL  FILL_223
timestamp 1018054153
transform 1 0 288 0 1 3140
box -16 -6 32 210
use FILL  FILL_224
timestamp 1018054153
transform 1 0 272 0 1 3140
box -16 -6 32 210
use FILL  FILL_225
timestamp 1018054153
transform 1 0 256 0 1 3140
box -16 -6 32 210
use FILL  FILL_226
timestamp 1018054153
transform 1 0 240 0 1 3140
box -16 -6 32 210
use FILL  FILL_227
timestamp 1018054153
transform 1 0 224 0 1 3140
box -16 -6 32 210
use FILL  FILL_228
timestamp 1018054153
transform 1 0 208 0 1 3140
box -16 -6 32 210
use FILL  FILL_229
timestamp 1018054153
transform 1 0 192 0 1 3140
box -16 -6 32 210
use FILL  FILL_230
timestamp 1018054153
transform 1 0 176 0 1 3140
box -16 -6 32 210
use FILL  FILL_231
timestamp 1018054153
transform 1 0 160 0 1 3140
box -16 -6 32 210
use FILL  FILL_232
timestamp 1018054153
transform 1 0 144 0 1 3140
box -16 -6 32 210
use FILL  FILL_233
timestamp 1018054153
transform 1 0 3664 0 -1 3140
box -16 -6 32 210
use FILL  FILL_234
timestamp 1018054153
transform 1 0 3648 0 -1 3140
box -16 -6 32 210
use FILL  FILL_235
timestamp 1018054153
transform 1 0 3632 0 -1 3140
box -16 -6 32 210
use FILL  FILL_236
timestamp 1018054153
transform 1 0 3616 0 -1 3140
box -16 -6 32 210
use FILL  FILL_237
timestamp 1018054153
transform 1 0 3600 0 -1 3140
box -16 -6 32 210
use FILL  FILL_238
timestamp 1018054153
transform 1 0 3584 0 -1 3140
box -16 -6 32 210
use FILL  FILL_239
timestamp 1018054153
transform 1 0 3568 0 -1 3140
box -16 -6 32 210
use FILL  FILL_240
timestamp 1018054153
transform 1 0 3552 0 -1 3140
box -16 -6 32 210
use FILL  FILL_241
timestamp 1018054153
transform 1 0 3536 0 -1 3140
box -16 -6 32 210
use FILL  FILL_242
timestamp 1018054153
transform 1 0 3520 0 -1 3140
box -16 -6 32 210
use FILL  FILL_243
timestamp 1018054153
transform 1 0 3504 0 -1 3140
box -16 -6 32 210
use FILL  FILL_244
timestamp 1018054153
transform 1 0 3488 0 -1 3140
box -16 -6 32 210
use FILL  FILL_245
timestamp 1018054153
transform 1 0 3472 0 -1 3140
box -16 -6 32 210
use FILL  FILL_246
timestamp 1018054153
transform 1 0 3456 0 -1 3140
box -16 -6 32 210
use FILL  FILL_247
timestamp 1018054153
transform 1 0 3440 0 -1 3140
box -16 -6 32 210
use FILL  FILL_248
timestamp 1018054153
transform 1 0 3424 0 -1 3140
box -16 -6 32 210
use FILL  FILL_249
timestamp 1018054153
transform 1 0 3408 0 -1 3140
box -16 -6 32 210
use FILL  FILL_250
timestamp 1018054153
transform 1 0 3392 0 -1 3140
box -16 -6 32 210
use FILL  FILL_251
timestamp 1018054153
transform 1 0 3376 0 -1 3140
box -16 -6 32 210
use FILL  FILL_252
timestamp 1018054153
transform 1 0 3360 0 -1 3140
box -16 -6 32 210
use FILL  FILL_253
timestamp 1018054153
transform 1 0 3344 0 -1 3140
box -16 -6 32 210
use FILL  FILL_254
timestamp 1018054153
transform 1 0 3328 0 -1 3140
box -16 -6 32 210
use FILL  FILL_255
timestamp 1018054153
transform 1 0 3312 0 -1 3140
box -16 -6 32 210
use FILL  FILL_256
timestamp 1018054153
transform 1 0 3264 0 -1 3140
box -16 -6 32 210
use FILL  FILL_257
timestamp 1018054153
transform 1 0 3248 0 -1 3140
box -16 -6 32 210
use FILL  FILL_258
timestamp 1018054153
transform 1 0 3152 0 -1 3140
box -16 -6 32 210
use FILL  FILL_259
timestamp 1018054153
transform 1 0 2640 0 -1 3140
box -16 -6 32 210
use FILL  FILL_260
timestamp 1018054153
transform 1 0 2080 0 -1 3140
box -16 -6 32 210
use FILL  FILL_261
timestamp 1018054153
transform 1 0 2064 0 -1 3140
box -16 -6 32 210
use FILL  FILL_262
timestamp 1018054153
transform 1 0 2048 0 -1 3140
box -16 -6 32 210
use FILL  FILL_263
timestamp 1018054153
transform 1 0 2032 0 -1 3140
box -16 -6 32 210
use FILL  FILL_264
timestamp 1018054153
transform 1 0 1952 0 -1 3140
box -16 -6 32 210
use FILL  FILL_265
timestamp 1018054153
transform 1 0 704 0 -1 3140
box -16 -6 32 210
use FILL  FILL_266
timestamp 1018054153
transform 1 0 688 0 -1 3140
box -16 -6 32 210
use FILL  FILL_267
timestamp 1018054153
transform 1 0 672 0 -1 3140
box -16 -6 32 210
use FILL  FILL_268
timestamp 1018054153
transform 1 0 656 0 -1 3140
box -16 -6 32 210
use FILL  FILL_269
timestamp 1018054153
transform 1 0 640 0 -1 3140
box -16 -6 32 210
use FILL  FILL_270
timestamp 1018054153
transform 1 0 624 0 -1 3140
box -16 -6 32 210
use FILL  FILL_271
timestamp 1018054153
transform 1 0 384 0 -1 3140
box -16 -6 32 210
use FILL  FILL_272
timestamp 1018054153
transform 1 0 336 0 -1 3140
box -16 -6 32 210
use FILL  FILL_273
timestamp 1018054153
transform 1 0 320 0 -1 3140
box -16 -6 32 210
use FILL  FILL_274
timestamp 1018054153
transform 1 0 304 0 -1 3140
box -16 -6 32 210
use FILL  FILL_275
timestamp 1018054153
transform 1 0 288 0 -1 3140
box -16 -6 32 210
use FILL  FILL_276
timestamp 1018054153
transform 1 0 272 0 -1 3140
box -16 -6 32 210
use FILL  FILL_277
timestamp 1018054153
transform 1 0 256 0 -1 3140
box -16 -6 32 210
use FILL  FILL_278
timestamp 1018054153
transform 1 0 240 0 -1 3140
box -16 -6 32 210
use FILL  FILL_279
timestamp 1018054153
transform 1 0 224 0 -1 3140
box -16 -6 32 210
use FILL  FILL_280
timestamp 1018054153
transform 1 0 208 0 -1 3140
box -16 -6 32 210
use FILL  FILL_281
timestamp 1018054153
transform 1 0 192 0 -1 3140
box -16 -6 32 210
use FILL  FILL_282
timestamp 1018054153
transform 1 0 176 0 -1 3140
box -16 -6 32 210
use FILL  FILL_283
timestamp 1018054153
transform 1 0 160 0 -1 3140
box -16 -6 32 210
use FILL  FILL_284
timestamp 1018054153
transform 1 0 144 0 -1 3140
box -16 -6 32 210
use FILL  FILL_285
timestamp 1018054153
transform 1 0 3664 0 1 2740
box -16 -6 32 210
use FILL  FILL_286
timestamp 1018054153
transform 1 0 3648 0 1 2740
box -16 -6 32 210
use FILL  FILL_287
timestamp 1018054153
transform 1 0 3632 0 1 2740
box -16 -6 32 210
use FILL  FILL_288
timestamp 1018054153
transform 1 0 3616 0 1 2740
box -16 -6 32 210
use FILL  FILL_289
timestamp 1018054153
transform 1 0 3600 0 1 2740
box -16 -6 32 210
use FILL  FILL_290
timestamp 1018054153
transform 1 0 3584 0 1 2740
box -16 -6 32 210
use FILL  FILL_291
timestamp 1018054153
transform 1 0 3568 0 1 2740
box -16 -6 32 210
use FILL  FILL_292
timestamp 1018054153
transform 1 0 3552 0 1 2740
box -16 -6 32 210
use FILL  FILL_293
timestamp 1018054153
transform 1 0 3536 0 1 2740
box -16 -6 32 210
use FILL  FILL_294
timestamp 1018054153
transform 1 0 3520 0 1 2740
box -16 -6 32 210
use FILL  FILL_295
timestamp 1018054153
transform 1 0 3504 0 1 2740
box -16 -6 32 210
use FILL  FILL_296
timestamp 1018054153
transform 1 0 3488 0 1 2740
box -16 -6 32 210
use FILL  FILL_297
timestamp 1018054153
transform 1 0 3472 0 1 2740
box -16 -6 32 210
use FILL  FILL_298
timestamp 1018054153
transform 1 0 3456 0 1 2740
box -16 -6 32 210
use FILL  FILL_299
timestamp 1018054153
transform 1 0 3440 0 1 2740
box -16 -6 32 210
use FILL  FILL_300
timestamp 1018054153
transform 1 0 3424 0 1 2740
box -16 -6 32 210
use FILL  FILL_301
timestamp 1018054153
transform 1 0 3408 0 1 2740
box -16 -6 32 210
use FILL  FILL_302
timestamp 1018054153
transform 1 0 3392 0 1 2740
box -16 -6 32 210
use FILL  FILL_303
timestamp 1018054153
transform 1 0 3376 0 1 2740
box -16 -6 32 210
use FILL  FILL_304
timestamp 1018054153
transform 1 0 3328 0 1 2740
box -16 -6 32 210
use FILL  FILL_305
timestamp 1018054153
transform 1 0 3232 0 1 2740
box -16 -6 32 210
use FILL  FILL_306
timestamp 1018054153
transform 1 0 3216 0 1 2740
box -16 -6 32 210
use FILL  FILL_307
timestamp 1018054153
transform 1 0 3200 0 1 2740
box -16 -6 32 210
use FILL  FILL_308
timestamp 1018054153
transform 1 0 3184 0 1 2740
box -16 -6 32 210
use FILL  FILL_309
timestamp 1018054153
transform 1 0 3168 0 1 2740
box -16 -6 32 210
use FILL  FILL_310
timestamp 1018054153
transform 1 0 3152 0 1 2740
box -16 -6 32 210
use FILL  FILL_311
timestamp 1018054153
transform 1 0 3136 0 1 2740
box -16 -6 32 210
use FILL  FILL_312
timestamp 1018054153
transform 1 0 1792 0 1 2740
box -16 -6 32 210
use FILL  FILL_313
timestamp 1018054153
transform 1 0 1712 0 1 2740
box -16 -6 32 210
use FILL  FILL_314
timestamp 1018054153
transform 1 0 1696 0 1 2740
box -16 -6 32 210
use FILL  FILL_315
timestamp 1018054153
transform 1 0 1680 0 1 2740
box -16 -6 32 210
use FILL  FILL_316
timestamp 1018054153
transform 1 0 1232 0 1 2740
box -16 -6 32 210
use FILL  FILL_317
timestamp 1018054153
transform 1 0 832 0 1 2740
box -16 -6 32 210
use FILL  FILL_318
timestamp 1018054153
transform 1 0 816 0 1 2740
box -16 -6 32 210
use FILL  FILL_319
timestamp 1018054153
transform 1 0 800 0 1 2740
box -16 -6 32 210
use FILL  FILL_320
timestamp 1018054153
transform 1 0 784 0 1 2740
box -16 -6 32 210
use FILL  FILL_321
timestamp 1018054153
transform 1 0 768 0 1 2740
box -16 -6 32 210
use FILL  FILL_322
timestamp 1018054153
transform 1 0 752 0 1 2740
box -16 -6 32 210
use FILL  FILL_323
timestamp 1018054153
transform 1 0 736 0 1 2740
box -16 -6 32 210
use FILL  FILL_324
timestamp 1018054153
transform 1 0 720 0 1 2740
box -16 -6 32 210
use FILL  FILL_325
timestamp 1018054153
transform 1 0 704 0 1 2740
box -16 -6 32 210
use FILL  FILL_326
timestamp 1018054153
transform 1 0 688 0 1 2740
box -16 -6 32 210
use FILL  FILL_327
timestamp 1018054153
transform 1 0 672 0 1 2740
box -16 -6 32 210
use FILL  FILL_328
timestamp 1018054153
transform 1 0 656 0 1 2740
box -16 -6 32 210
use FILL  FILL_329
timestamp 1018054153
transform 1 0 496 0 1 2740
box -16 -6 32 210
use FILL  FILL_330
timestamp 1018054153
transform 1 0 480 0 1 2740
box -16 -6 32 210
use FILL  FILL_331
timestamp 1018054153
transform 1 0 464 0 1 2740
box -16 -6 32 210
use FILL  FILL_332
timestamp 1018054153
transform 1 0 448 0 1 2740
box -16 -6 32 210
use FILL  FILL_333
timestamp 1018054153
transform 1 0 432 0 1 2740
box -16 -6 32 210
use FILL  FILL_334
timestamp 1018054153
transform 1 0 416 0 1 2740
box -16 -6 32 210
use FILL  FILL_335
timestamp 1018054153
transform 1 0 400 0 1 2740
box -16 -6 32 210
use FILL  FILL_336
timestamp 1018054153
transform 1 0 384 0 1 2740
box -16 -6 32 210
use FILL  FILL_337
timestamp 1018054153
transform 1 0 368 0 1 2740
box -16 -6 32 210
use FILL  FILL_338
timestamp 1018054153
transform 1 0 352 0 1 2740
box -16 -6 32 210
use FILL  FILL_339
timestamp 1018054153
transform 1 0 336 0 1 2740
box -16 -6 32 210
use FILL  FILL_340
timestamp 1018054153
transform 1 0 320 0 1 2740
box -16 -6 32 210
use FILL  FILL_341
timestamp 1018054153
transform 1 0 304 0 1 2740
box -16 -6 32 210
use FILL  FILL_342
timestamp 1018054153
transform 1 0 288 0 1 2740
box -16 -6 32 210
use FILL  FILL_343
timestamp 1018054153
transform 1 0 272 0 1 2740
box -16 -6 32 210
use FILL  FILL_344
timestamp 1018054153
transform 1 0 256 0 1 2740
box -16 -6 32 210
use FILL  FILL_345
timestamp 1018054153
transform 1 0 240 0 1 2740
box -16 -6 32 210
use FILL  FILL_346
timestamp 1018054153
transform 1 0 224 0 1 2740
box -16 -6 32 210
use FILL  FILL_347
timestamp 1018054153
transform 1 0 208 0 1 2740
box -16 -6 32 210
use FILL  FILL_348
timestamp 1018054153
transform 1 0 192 0 1 2740
box -16 -6 32 210
use FILL  FILL_349
timestamp 1018054153
transform 1 0 176 0 1 2740
box -16 -6 32 210
use FILL  FILL_350
timestamp 1018054153
transform 1 0 160 0 1 2740
box -16 -6 32 210
use FILL  FILL_351
timestamp 1018054153
transform 1 0 144 0 1 2740
box -16 -6 32 210
use FILL  FILL_352
timestamp 1018054153
transform 1 0 3664 0 -1 2740
box -16 -6 32 210
use FILL  FILL_353
timestamp 1018054153
transform 1 0 3648 0 -1 2740
box -16 -6 32 210
use FILL  FILL_354
timestamp 1018054153
transform 1 0 3632 0 -1 2740
box -16 -6 32 210
use FILL  FILL_355
timestamp 1018054153
transform 1 0 3616 0 -1 2740
box -16 -6 32 210
use FILL  FILL_356
timestamp 1018054153
transform 1 0 3600 0 -1 2740
box -16 -6 32 210
use FILL  FILL_357
timestamp 1018054153
transform 1 0 3584 0 -1 2740
box -16 -6 32 210
use FILL  FILL_358
timestamp 1018054153
transform 1 0 3568 0 -1 2740
box -16 -6 32 210
use FILL  FILL_359
timestamp 1018054153
transform 1 0 3552 0 -1 2740
box -16 -6 32 210
use FILL  FILL_360
timestamp 1018054153
transform 1 0 3536 0 -1 2740
box -16 -6 32 210
use FILL  FILL_361
timestamp 1018054153
transform 1 0 3520 0 -1 2740
box -16 -6 32 210
use FILL  FILL_362
timestamp 1018054153
transform 1 0 3504 0 -1 2740
box -16 -6 32 210
use FILL  FILL_363
timestamp 1018054153
transform 1 0 3488 0 -1 2740
box -16 -6 32 210
use FILL  FILL_364
timestamp 1018054153
transform 1 0 3472 0 -1 2740
box -16 -6 32 210
use FILL  FILL_365
timestamp 1018054153
transform 1 0 3456 0 -1 2740
box -16 -6 32 210
use FILL  FILL_366
timestamp 1018054153
transform 1 0 3440 0 -1 2740
box -16 -6 32 210
use FILL  FILL_367
timestamp 1018054153
transform 1 0 3424 0 -1 2740
box -16 -6 32 210
use FILL  FILL_368
timestamp 1018054153
transform 1 0 3408 0 -1 2740
box -16 -6 32 210
use FILL  FILL_369
timestamp 1018054153
transform 1 0 3392 0 -1 2740
box -16 -6 32 210
use FILL  FILL_370
timestamp 1018054153
transform 1 0 3376 0 -1 2740
box -16 -6 32 210
use FILL  FILL_371
timestamp 1018054153
transform 1 0 3360 0 -1 2740
box -16 -6 32 210
use FILL  FILL_372
timestamp 1018054153
transform 1 0 1920 0 -1 2740
box -16 -6 32 210
use FILL  FILL_373
timestamp 1018054153
transform 1 0 1904 0 -1 2740
box -16 -6 32 210
use FILL  FILL_374
timestamp 1018054153
transform 1 0 1808 0 -1 2740
box -16 -6 32 210
use FILL  FILL_375
timestamp 1018054153
transform 1 0 576 0 -1 2740
box -16 -6 32 210
use FILL  FILL_376
timestamp 1018054153
transform 1 0 560 0 -1 2740
box -16 -6 32 210
use FILL  FILL_377
timestamp 1018054153
transform 1 0 512 0 -1 2740
box -16 -6 32 210
use FILL  FILL_378
timestamp 1018054153
transform 1 0 496 0 -1 2740
box -16 -6 32 210
use FILL  FILL_379
timestamp 1018054153
transform 1 0 480 0 -1 2740
box -16 -6 32 210
use FILL  FILL_380
timestamp 1018054153
transform 1 0 464 0 -1 2740
box -16 -6 32 210
use FILL  FILL_381
timestamp 1018054153
transform 1 0 448 0 -1 2740
box -16 -6 32 210
use FILL  FILL_382
timestamp 1018054153
transform 1 0 432 0 -1 2740
box -16 -6 32 210
use FILL  FILL_383
timestamp 1018054153
transform 1 0 416 0 -1 2740
box -16 -6 32 210
use FILL  FILL_384
timestamp 1018054153
transform 1 0 400 0 -1 2740
box -16 -6 32 210
use FILL  FILL_385
timestamp 1018054153
transform 1 0 384 0 -1 2740
box -16 -6 32 210
use FILL  FILL_386
timestamp 1018054153
transform 1 0 368 0 -1 2740
box -16 -6 32 210
use FILL  FILL_387
timestamp 1018054153
transform 1 0 352 0 -1 2740
box -16 -6 32 210
use FILL  FILL_388
timestamp 1018054153
transform 1 0 336 0 -1 2740
box -16 -6 32 210
use FILL  FILL_389
timestamp 1018054153
transform 1 0 320 0 -1 2740
box -16 -6 32 210
use FILL  FILL_390
timestamp 1018054153
transform 1 0 304 0 -1 2740
box -16 -6 32 210
use FILL  FILL_391
timestamp 1018054153
transform 1 0 288 0 -1 2740
box -16 -6 32 210
use FILL  FILL_392
timestamp 1018054153
transform 1 0 272 0 -1 2740
box -16 -6 32 210
use FILL  FILL_393
timestamp 1018054153
transform 1 0 256 0 -1 2740
box -16 -6 32 210
use FILL  FILL_394
timestamp 1018054153
transform 1 0 240 0 -1 2740
box -16 -6 32 210
use FILL  FILL_395
timestamp 1018054153
transform 1 0 224 0 -1 2740
box -16 -6 32 210
use FILL  FILL_396
timestamp 1018054153
transform 1 0 208 0 -1 2740
box -16 -6 32 210
use FILL  FILL_397
timestamp 1018054153
transform 1 0 192 0 -1 2740
box -16 -6 32 210
use FILL  FILL_398
timestamp 1018054153
transform 1 0 176 0 -1 2740
box -16 -6 32 210
use FILL  FILL_399
timestamp 1018054153
transform 1 0 160 0 -1 2740
box -16 -6 32 210
use FILL  FILL_400
timestamp 1018054153
transform 1 0 144 0 -1 2740
box -16 -6 32 210
use FILL  FILL_401
timestamp 1018054153
transform 1 0 3664 0 1 2340
box -16 -6 32 210
use FILL  FILL_402
timestamp 1018054153
transform 1 0 3648 0 1 2340
box -16 -6 32 210
use FILL  FILL_403
timestamp 1018054153
transform 1 0 3632 0 1 2340
box -16 -6 32 210
use FILL  FILL_404
timestamp 1018054153
transform 1 0 3616 0 1 2340
box -16 -6 32 210
use FILL  FILL_405
timestamp 1018054153
transform 1 0 3600 0 1 2340
box -16 -6 32 210
use FILL  FILL_406
timestamp 1018054153
transform 1 0 3584 0 1 2340
box -16 -6 32 210
use FILL  FILL_407
timestamp 1018054153
transform 1 0 3568 0 1 2340
box -16 -6 32 210
use FILL  FILL_408
timestamp 1018054153
transform 1 0 3552 0 1 2340
box -16 -6 32 210
use FILL  FILL_409
timestamp 1018054153
transform 1 0 3536 0 1 2340
box -16 -6 32 210
use FILL  FILL_410
timestamp 1018054153
transform 1 0 3520 0 1 2340
box -16 -6 32 210
use FILL  FILL_411
timestamp 1018054153
transform 1 0 3504 0 1 2340
box -16 -6 32 210
use FILL  FILL_412
timestamp 1018054153
transform 1 0 3488 0 1 2340
box -16 -6 32 210
use FILL  FILL_413
timestamp 1018054153
transform 1 0 3472 0 1 2340
box -16 -6 32 210
use FILL  FILL_414
timestamp 1018054153
transform 1 0 3456 0 1 2340
box -16 -6 32 210
use FILL  FILL_415
timestamp 1018054153
transform 1 0 3440 0 1 2340
box -16 -6 32 210
use FILL  FILL_416
timestamp 1018054153
transform 1 0 3424 0 1 2340
box -16 -6 32 210
use FILL  FILL_417
timestamp 1018054153
transform 1 0 3408 0 1 2340
box -16 -6 32 210
use FILL  FILL_418
timestamp 1018054153
transform 1 0 3392 0 1 2340
box -16 -6 32 210
use FILL  FILL_419
timestamp 1018054153
transform 1 0 3376 0 1 2340
box -16 -6 32 210
use FILL  FILL_420
timestamp 1018054153
transform 1 0 3360 0 1 2340
box -16 -6 32 210
use FILL  FILL_421
timestamp 1018054153
transform 1 0 3344 0 1 2340
box -16 -6 32 210
use FILL  FILL_422
timestamp 1018054153
transform 1 0 3328 0 1 2340
box -16 -6 32 210
use FILL  FILL_423
timestamp 1018054153
transform 1 0 3312 0 1 2340
box -16 -6 32 210
use FILL  FILL_424
timestamp 1018054153
transform 1 0 3296 0 1 2340
box -16 -6 32 210
use FILL  FILL_425
timestamp 1018054153
transform 1 0 3280 0 1 2340
box -16 -6 32 210
use FILL  FILL_426
timestamp 1018054153
transform 1 0 3264 0 1 2340
box -16 -6 32 210
use FILL  FILL_427
timestamp 1018054153
transform 1 0 3248 0 1 2340
box -16 -6 32 210
use FILL  FILL_428
timestamp 1018054153
transform 1 0 3232 0 1 2340
box -16 -6 32 210
use FILL  FILL_429
timestamp 1018054153
transform 1 0 3216 0 1 2340
box -16 -6 32 210
use FILL  FILL_430
timestamp 1018054153
transform 1 0 3200 0 1 2340
box -16 -6 32 210
use FILL  FILL_431
timestamp 1018054153
transform 1 0 3184 0 1 2340
box -16 -6 32 210
use FILL  FILL_432
timestamp 1018054153
transform 1 0 3168 0 1 2340
box -16 -6 32 210
use FILL  FILL_433
timestamp 1018054153
transform 1 0 3152 0 1 2340
box -16 -6 32 210
use FILL  FILL_434
timestamp 1018054153
transform 1 0 3136 0 1 2340
box -16 -6 32 210
use FILL  FILL_435
timestamp 1018054153
transform 1 0 3120 0 1 2340
box -16 -6 32 210
use FILL  FILL_436
timestamp 1018054153
transform 1 0 3104 0 1 2340
box -16 -6 32 210
use FILL  FILL_437
timestamp 1018054153
transform 1 0 2976 0 1 2340
box -16 -6 32 210
use FILL  FILL_438
timestamp 1018054153
transform 1 0 2960 0 1 2340
box -16 -6 32 210
use FILL  FILL_439
timestamp 1018054153
transform 1 0 2944 0 1 2340
box -16 -6 32 210
use FILL  FILL_440
timestamp 1018054153
transform 1 0 2928 0 1 2340
box -16 -6 32 210
use FILL  FILL_441
timestamp 1018054153
transform 1 0 2912 0 1 2340
box -16 -6 32 210
use FILL  FILL_442
timestamp 1018054153
transform 1 0 2896 0 1 2340
box -16 -6 32 210
use FILL  FILL_443
timestamp 1018054153
transform 1 0 2880 0 1 2340
box -16 -6 32 210
use FILL  FILL_444
timestamp 1018054153
transform 1 0 2704 0 1 2340
box -16 -6 32 210
use FILL  FILL_445
timestamp 1018054153
transform 1 0 2688 0 1 2340
box -16 -6 32 210
use FILL  FILL_446
timestamp 1018054153
transform 1 0 2672 0 1 2340
box -16 -6 32 210
use FILL  FILL_447
timestamp 1018054153
transform 1 0 2384 0 1 2340
box -16 -6 32 210
use FILL  FILL_448
timestamp 1018054153
transform 1 0 2096 0 1 2340
box -16 -6 32 210
use FILL  FILL_449
timestamp 1018054153
transform 1 0 2080 0 1 2340
box -16 -6 32 210
use FILL  FILL_450
timestamp 1018054153
transform 1 0 2064 0 1 2340
box -16 -6 32 210
use FILL  FILL_451
timestamp 1018054153
transform 1 0 2048 0 1 2340
box -16 -6 32 210
use FILL  FILL_452
timestamp 1018054153
transform 1 0 1952 0 1 2340
box -16 -6 32 210
use FILL  FILL_453
timestamp 1018054153
transform 1 0 1936 0 1 2340
box -16 -6 32 210
use FILL  FILL_454
timestamp 1018054153
transform 1 0 1920 0 1 2340
box -16 -6 32 210
use FILL  FILL_455
timestamp 1018054153
transform 1 0 1904 0 1 2340
box -16 -6 32 210
use FILL  FILL_456
timestamp 1018054153
transform 1 0 1808 0 1 2340
box -16 -6 32 210
use FILL  FILL_457
timestamp 1018054153
transform 1 0 1792 0 1 2340
box -16 -6 32 210
use FILL  FILL_458
timestamp 1018054153
transform 1 0 1776 0 1 2340
box -16 -6 32 210
use FILL  FILL_459
timestamp 1018054153
transform 1 0 1760 0 1 2340
box -16 -6 32 210
use FILL  FILL_460
timestamp 1018054153
transform 1 0 1744 0 1 2340
box -16 -6 32 210
use FILL  FILL_461
timestamp 1018054153
transform 1 0 1728 0 1 2340
box -16 -6 32 210
use FILL  FILL_462
timestamp 1018054153
transform 1 0 1712 0 1 2340
box -16 -6 32 210
use FILL  FILL_463
timestamp 1018054153
transform 1 0 1536 0 1 2340
box -16 -6 32 210
use FILL  FILL_464
timestamp 1018054153
transform 1 0 1520 0 1 2340
box -16 -6 32 210
use FILL  FILL_465
timestamp 1018054153
transform 1 0 1504 0 1 2340
box -16 -6 32 210
use FILL  FILL_466
timestamp 1018054153
transform 1 0 1488 0 1 2340
box -16 -6 32 210
use FILL  FILL_467
timestamp 1018054153
transform 1 0 1312 0 1 2340
box -16 -6 32 210
use FILL  FILL_468
timestamp 1018054153
transform 1 0 1184 0 1 2340
box -16 -6 32 210
use FILL  FILL_469
timestamp 1018054153
transform 1 0 1168 0 1 2340
box -16 -6 32 210
use FILL  FILL_470
timestamp 1018054153
transform 1 0 1152 0 1 2340
box -16 -6 32 210
use FILL  FILL_471
timestamp 1018054153
transform 1 0 992 0 1 2340
box -16 -6 32 210
use FILL  FILL_472
timestamp 1018054153
transform 1 0 976 0 1 2340
box -16 -6 32 210
use FILL  FILL_473
timestamp 1018054153
transform 1 0 768 0 1 2340
box -16 -6 32 210
use FILL  FILL_474
timestamp 1018054153
transform 1 0 752 0 1 2340
box -16 -6 32 210
use FILL  FILL_475
timestamp 1018054153
transform 1 0 656 0 1 2340
box -16 -6 32 210
use FILL  FILL_476
timestamp 1018054153
transform 1 0 640 0 1 2340
box -16 -6 32 210
use FILL  FILL_477
timestamp 1018054153
transform 1 0 624 0 1 2340
box -16 -6 32 210
use FILL  FILL_478
timestamp 1018054153
transform 1 0 608 0 1 2340
box -16 -6 32 210
use FILL  FILL_479
timestamp 1018054153
transform 1 0 560 0 1 2340
box -16 -6 32 210
use FILL  FILL_480
timestamp 1018054153
transform 1 0 544 0 1 2340
box -16 -6 32 210
use FILL  FILL_481
timestamp 1018054153
transform 1 0 528 0 1 2340
box -16 -6 32 210
use FILL  FILL_482
timestamp 1018054153
transform 1 0 512 0 1 2340
box -16 -6 32 210
use FILL  FILL_483
timestamp 1018054153
transform 1 0 496 0 1 2340
box -16 -6 32 210
use FILL  FILL_484
timestamp 1018054153
transform 1 0 480 0 1 2340
box -16 -6 32 210
use FILL  FILL_485
timestamp 1018054153
transform 1 0 464 0 1 2340
box -16 -6 32 210
use FILL  FILL_486
timestamp 1018054153
transform 1 0 448 0 1 2340
box -16 -6 32 210
use FILL  FILL_487
timestamp 1018054153
transform 1 0 432 0 1 2340
box -16 -6 32 210
use FILL  FILL_488
timestamp 1018054153
transform 1 0 416 0 1 2340
box -16 -6 32 210
use FILL  FILL_489
timestamp 1018054153
transform 1 0 400 0 1 2340
box -16 -6 32 210
use FILL  FILL_490
timestamp 1018054153
transform 1 0 384 0 1 2340
box -16 -6 32 210
use FILL  FILL_491
timestamp 1018054153
transform 1 0 368 0 1 2340
box -16 -6 32 210
use FILL  FILL_492
timestamp 1018054153
transform 1 0 352 0 1 2340
box -16 -6 32 210
use FILL  FILL_493
timestamp 1018054153
transform 1 0 336 0 1 2340
box -16 -6 32 210
use FILL  FILL_494
timestamp 1018054153
transform 1 0 320 0 1 2340
box -16 -6 32 210
use FILL  FILL_495
timestamp 1018054153
transform 1 0 304 0 1 2340
box -16 -6 32 210
use FILL  FILL_496
timestamp 1018054153
transform 1 0 288 0 1 2340
box -16 -6 32 210
use FILL  FILL_497
timestamp 1018054153
transform 1 0 272 0 1 2340
box -16 -6 32 210
use FILL  FILL_498
timestamp 1018054153
transform 1 0 256 0 1 2340
box -16 -6 32 210
use FILL  FILL_499
timestamp 1018054153
transform 1 0 240 0 1 2340
box -16 -6 32 210
use FILL  FILL_500
timestamp 1018054153
transform 1 0 224 0 1 2340
box -16 -6 32 210
use FILL  FILL_501
timestamp 1018054153
transform 1 0 208 0 1 2340
box -16 -6 32 210
use FILL  FILL_502
timestamp 1018054153
transform 1 0 192 0 1 2340
box -16 -6 32 210
use FILL  FILL_503
timestamp 1018054153
transform 1 0 176 0 1 2340
box -16 -6 32 210
use FILL  FILL_504
timestamp 1018054153
transform 1 0 160 0 1 2340
box -16 -6 32 210
use FILL  FILL_505
timestamp 1018054153
transform 1 0 144 0 1 2340
box -16 -6 32 210
use FILL  FILL_506
timestamp 1018054153
transform 1 0 3664 0 -1 2340
box -16 -6 32 210
use FILL  FILL_507
timestamp 1018054153
transform 1 0 3648 0 -1 2340
box -16 -6 32 210
use FILL  FILL_508
timestamp 1018054153
transform 1 0 3632 0 -1 2340
box -16 -6 32 210
use FILL  FILL_509
timestamp 1018054153
transform 1 0 3616 0 -1 2340
box -16 -6 32 210
use FILL  FILL_510
timestamp 1018054153
transform 1 0 3600 0 -1 2340
box -16 -6 32 210
use FILL  FILL_511
timestamp 1018054153
transform 1 0 3584 0 -1 2340
box -16 -6 32 210
use FILL  FILL_512
timestamp 1018054153
transform 1 0 3568 0 -1 2340
box -16 -6 32 210
use FILL  FILL_513
timestamp 1018054153
transform 1 0 3552 0 -1 2340
box -16 -6 32 210
use FILL  FILL_514
timestamp 1018054153
transform 1 0 3536 0 -1 2340
box -16 -6 32 210
use FILL  FILL_515
timestamp 1018054153
transform 1 0 3520 0 -1 2340
box -16 -6 32 210
use FILL  FILL_516
timestamp 1018054153
transform 1 0 3504 0 -1 2340
box -16 -6 32 210
use FILL  FILL_517
timestamp 1018054153
transform 1 0 3488 0 -1 2340
box -16 -6 32 210
use FILL  FILL_518
timestamp 1018054153
transform 1 0 3472 0 -1 2340
box -16 -6 32 210
use FILL  FILL_519
timestamp 1018054153
transform 1 0 3456 0 -1 2340
box -16 -6 32 210
use FILL  FILL_520
timestamp 1018054153
transform 1 0 3440 0 -1 2340
box -16 -6 32 210
use FILL  FILL_521
timestamp 1018054153
transform 1 0 3424 0 -1 2340
box -16 -6 32 210
use FILL  FILL_522
timestamp 1018054153
transform 1 0 3408 0 -1 2340
box -16 -6 32 210
use FILL  FILL_523
timestamp 1018054153
transform 1 0 3392 0 -1 2340
box -16 -6 32 210
use FILL  FILL_524
timestamp 1018054153
transform 1 0 3376 0 -1 2340
box -16 -6 32 210
use FILL  FILL_525
timestamp 1018054153
transform 1 0 3360 0 -1 2340
box -16 -6 32 210
use FILL  FILL_526
timestamp 1018054153
transform 1 0 3344 0 -1 2340
box -16 -6 32 210
use FILL  FILL_527
timestamp 1018054153
transform 1 0 3328 0 -1 2340
box -16 -6 32 210
use FILL  FILL_528
timestamp 1018054153
transform 1 0 3312 0 -1 2340
box -16 -6 32 210
use FILL  FILL_529
timestamp 1018054153
transform 1 0 3296 0 -1 2340
box -16 -6 32 210
use FILL  FILL_530
timestamp 1018054153
transform 1 0 3280 0 -1 2340
box -16 -6 32 210
use FILL  FILL_531
timestamp 1018054153
transform 1 0 3040 0 -1 2340
box -16 -6 32 210
use FILL  FILL_532
timestamp 1018054153
transform 1 0 3024 0 -1 2340
box -16 -6 32 210
use FILL  FILL_533
timestamp 1018054153
transform 1 0 2896 0 -1 2340
box -16 -6 32 210
use FILL  FILL_534
timestamp 1018054153
transform 1 0 2880 0 -1 2340
box -16 -6 32 210
use FILL  FILL_535
timestamp 1018054153
transform 1 0 2864 0 -1 2340
box -16 -6 32 210
use FILL  FILL_536
timestamp 1018054153
transform 1 0 2848 0 -1 2340
box -16 -6 32 210
use FILL  FILL_537
timestamp 1018054153
transform 1 0 2832 0 -1 2340
box -16 -6 32 210
use FILL  FILL_538
timestamp 1018054153
transform 1 0 2816 0 -1 2340
box -16 -6 32 210
use FILL  FILL_539
timestamp 1018054153
transform 1 0 2688 0 -1 2340
box -16 -6 32 210
use FILL  FILL_540
timestamp 1018054153
transform 1 0 2672 0 -1 2340
box -16 -6 32 210
use FILL  FILL_541
timestamp 1018054153
transform 1 0 2656 0 -1 2340
box -16 -6 32 210
use FILL  FILL_542
timestamp 1018054153
transform 1 0 2640 0 -1 2340
box -16 -6 32 210
use FILL  FILL_543
timestamp 1018054153
transform 1 0 2624 0 -1 2340
box -16 -6 32 210
use FILL  FILL_544
timestamp 1018054153
transform 1 0 2496 0 -1 2340
box -16 -6 32 210
use FILL  FILL_545
timestamp 1018054153
transform 1 0 2480 0 -1 2340
box -16 -6 32 210
use FILL  FILL_546
timestamp 1018054153
transform 1 0 2304 0 -1 2340
box -16 -6 32 210
use FILL  FILL_547
timestamp 1018054153
transform 1 0 2288 0 -1 2340
box -16 -6 32 210
use FILL  FILL_548
timestamp 1018054153
transform 1 0 2272 0 -1 2340
box -16 -6 32 210
use FILL  FILL_549
timestamp 1018054153
transform 1 0 2256 0 -1 2340
box -16 -6 32 210
use FILL  FILL_550
timestamp 1018054153
transform 1 0 2240 0 -1 2340
box -16 -6 32 210
use FILL  FILL_551
timestamp 1018054153
transform 1 0 2224 0 -1 2340
box -16 -6 32 210
use FILL  FILL_552
timestamp 1018054153
transform 1 0 2208 0 -1 2340
box -16 -6 32 210
use FILL  FILL_553
timestamp 1018054153
transform 1 0 2192 0 -1 2340
box -16 -6 32 210
use FILL  FILL_554
timestamp 1018054153
transform 1 0 2176 0 -1 2340
box -16 -6 32 210
use FILL  FILL_555
timestamp 1018054153
transform 1 0 2160 0 -1 2340
box -16 -6 32 210
use FILL  FILL_556
timestamp 1018054153
transform 1 0 1920 0 -1 2340
box -16 -6 32 210
use FILL  FILL_557
timestamp 1018054153
transform 1 0 1904 0 -1 2340
box -16 -6 32 210
use FILL  FILL_558
timestamp 1018054153
transform 1 0 1616 0 -1 2340
box -16 -6 32 210
use FILL  FILL_559
timestamp 1018054153
transform 1 0 1600 0 -1 2340
box -16 -6 32 210
use FILL  FILL_560
timestamp 1018054153
transform 1 0 1584 0 -1 2340
box -16 -6 32 210
use FILL  FILL_561
timestamp 1018054153
transform 1 0 1408 0 -1 2340
box -16 -6 32 210
use FILL  FILL_562
timestamp 1018054153
transform 1 0 1280 0 -1 2340
box -16 -6 32 210
use FILL  FILL_563
timestamp 1018054153
transform 1 0 1264 0 -1 2340
box -16 -6 32 210
use FILL  FILL_564
timestamp 1018054153
transform 1 0 1248 0 -1 2340
box -16 -6 32 210
use FILL  FILL_565
timestamp 1018054153
transform 1 0 1088 0 -1 2340
box -16 -6 32 210
use FILL  FILL_566
timestamp 1018054153
transform 1 0 1072 0 -1 2340
box -16 -6 32 210
use FILL  FILL_567
timestamp 1018054153
transform 1 0 1056 0 -1 2340
box -16 -6 32 210
use FILL  FILL_568
timestamp 1018054153
transform 1 0 864 0 -1 2340
box -16 -6 32 210
use FILL  FILL_569
timestamp 1018054153
transform 1 0 848 0 -1 2340
box -16 -6 32 210
use FILL  FILL_570
timestamp 1018054153
transform 1 0 832 0 -1 2340
box -16 -6 32 210
use FILL  FILL_571
timestamp 1018054153
transform 1 0 816 0 -1 2340
box -16 -6 32 210
use FILL  FILL_572
timestamp 1018054153
transform 1 0 576 0 -1 2340
box -16 -6 32 210
use FILL  FILL_573
timestamp 1018054153
transform 1 0 560 0 -1 2340
box -16 -6 32 210
use FILL  FILL_574
timestamp 1018054153
transform 1 0 544 0 -1 2340
box -16 -6 32 210
use FILL  FILL_575
timestamp 1018054153
transform 1 0 528 0 -1 2340
box -16 -6 32 210
use FILL  FILL_576
timestamp 1018054153
transform 1 0 512 0 -1 2340
box -16 -6 32 210
use FILL  FILL_577
timestamp 1018054153
transform 1 0 496 0 -1 2340
box -16 -6 32 210
use FILL  FILL_578
timestamp 1018054153
transform 1 0 480 0 -1 2340
box -16 -6 32 210
use FILL  FILL_579
timestamp 1018054153
transform 1 0 464 0 -1 2340
box -16 -6 32 210
use FILL  FILL_580
timestamp 1018054153
transform 1 0 448 0 -1 2340
box -16 -6 32 210
use FILL  FILL_581
timestamp 1018054153
transform 1 0 432 0 -1 2340
box -16 -6 32 210
use FILL  FILL_582
timestamp 1018054153
transform 1 0 416 0 -1 2340
box -16 -6 32 210
use FILL  FILL_583
timestamp 1018054153
transform 1 0 400 0 -1 2340
box -16 -6 32 210
use FILL  FILL_584
timestamp 1018054153
transform 1 0 384 0 -1 2340
box -16 -6 32 210
use FILL  FILL_585
timestamp 1018054153
transform 1 0 368 0 -1 2340
box -16 -6 32 210
use FILL  FILL_586
timestamp 1018054153
transform 1 0 352 0 -1 2340
box -16 -6 32 210
use FILL  FILL_587
timestamp 1018054153
transform 1 0 336 0 -1 2340
box -16 -6 32 210
use FILL  FILL_588
timestamp 1018054153
transform 1 0 320 0 -1 2340
box -16 -6 32 210
use FILL  FILL_589
timestamp 1018054153
transform 1 0 304 0 -1 2340
box -16 -6 32 210
use FILL  FILL_590
timestamp 1018054153
transform 1 0 288 0 -1 2340
box -16 -6 32 210
use FILL  FILL_591
timestamp 1018054153
transform 1 0 272 0 -1 2340
box -16 -6 32 210
use FILL  FILL_592
timestamp 1018054153
transform 1 0 256 0 -1 2340
box -16 -6 32 210
use FILL  FILL_593
timestamp 1018054153
transform 1 0 240 0 -1 2340
box -16 -6 32 210
use FILL  FILL_594
timestamp 1018054153
transform 1 0 224 0 -1 2340
box -16 -6 32 210
use FILL  FILL_595
timestamp 1018054153
transform 1 0 208 0 -1 2340
box -16 -6 32 210
use FILL  FILL_596
timestamp 1018054153
transform 1 0 192 0 -1 2340
box -16 -6 32 210
use FILL  FILL_597
timestamp 1018054153
transform 1 0 176 0 -1 2340
box -16 -6 32 210
use FILL  FILL_598
timestamp 1018054153
transform 1 0 160 0 -1 2340
box -16 -6 32 210
use FILL  FILL_599
timestamp 1018054153
transform 1 0 144 0 -1 2340
box -16 -6 32 210
use FILL  FILL_600
timestamp 1018054153
transform 1 0 3664 0 1 1940
box -16 -6 32 210
use FILL  FILL_601
timestamp 1018054153
transform 1 0 3648 0 1 1940
box -16 -6 32 210
use FILL  FILL_602
timestamp 1018054153
transform 1 0 3632 0 1 1940
box -16 -6 32 210
use FILL  FILL_603
timestamp 1018054153
transform 1 0 3616 0 1 1940
box -16 -6 32 210
use FILL  FILL_604
timestamp 1018054153
transform 1 0 3600 0 1 1940
box -16 -6 32 210
use FILL  FILL_605
timestamp 1018054153
transform 1 0 3584 0 1 1940
box -16 -6 32 210
use FILL  FILL_606
timestamp 1018054153
transform 1 0 3568 0 1 1940
box -16 -6 32 210
use FILL  FILL_607
timestamp 1018054153
transform 1 0 3552 0 1 1940
box -16 -6 32 210
use FILL  FILL_608
timestamp 1018054153
transform 1 0 3536 0 1 1940
box -16 -6 32 210
use FILL  FILL_609
timestamp 1018054153
transform 1 0 3520 0 1 1940
box -16 -6 32 210
use FILL  FILL_610
timestamp 1018054153
transform 1 0 3504 0 1 1940
box -16 -6 32 210
use FILL  FILL_611
timestamp 1018054153
transform 1 0 3488 0 1 1940
box -16 -6 32 210
use FILL  FILL_612
timestamp 1018054153
transform 1 0 3472 0 1 1940
box -16 -6 32 210
use FILL  FILL_613
timestamp 1018054153
transform 1 0 3456 0 1 1940
box -16 -6 32 210
use FILL  FILL_614
timestamp 1018054153
transform 1 0 3440 0 1 1940
box -16 -6 32 210
use FILL  FILL_615
timestamp 1018054153
transform 1 0 3424 0 1 1940
box -16 -6 32 210
use FILL  FILL_616
timestamp 1018054153
transform 1 0 3408 0 1 1940
box -16 -6 32 210
use FILL  FILL_617
timestamp 1018054153
transform 1 0 3392 0 1 1940
box -16 -6 32 210
use FILL  FILL_618
timestamp 1018054153
transform 1 0 3376 0 1 1940
box -16 -6 32 210
use FILL  FILL_619
timestamp 1018054153
transform 1 0 3360 0 1 1940
box -16 -6 32 210
use FILL  FILL_620
timestamp 1018054153
transform 1 0 3344 0 1 1940
box -16 -6 32 210
use FILL  FILL_621
timestamp 1018054153
transform 1 0 3328 0 1 1940
box -16 -6 32 210
use FILL  FILL_622
timestamp 1018054153
transform 1 0 3312 0 1 1940
box -16 -6 32 210
use FILL  FILL_623
timestamp 1018054153
transform 1 0 3296 0 1 1940
box -16 -6 32 210
use FILL  FILL_624
timestamp 1018054153
transform 1 0 3280 0 1 1940
box -16 -6 32 210
use FILL  FILL_625
timestamp 1018054153
transform 1 0 3184 0 1 1940
box -16 -6 32 210
use FILL  FILL_626
timestamp 1018054153
transform 1 0 3168 0 1 1940
box -16 -6 32 210
use FILL  FILL_627
timestamp 1018054153
transform 1 0 3152 0 1 1940
box -16 -6 32 210
use FILL  FILL_628
timestamp 1018054153
transform 1 0 3136 0 1 1940
box -16 -6 32 210
use FILL  FILL_629
timestamp 1018054153
transform 1 0 3120 0 1 1940
box -16 -6 32 210
use FILL  FILL_630
timestamp 1018054153
transform 1 0 3104 0 1 1940
box -16 -6 32 210
use FILL  FILL_631
timestamp 1018054153
transform 1 0 3088 0 1 1940
box -16 -6 32 210
use FILL  FILL_632
timestamp 1018054153
transform 1 0 3072 0 1 1940
box -16 -6 32 210
use FILL  FILL_633
timestamp 1018054153
transform 1 0 3024 0 1 1940
box -16 -6 32 210
use FILL  FILL_634
timestamp 1018054153
transform 1 0 3008 0 1 1940
box -16 -6 32 210
use FILL  FILL_635
timestamp 1018054153
transform 1 0 2912 0 1 1940
box -16 -6 32 210
use FILL  FILL_636
timestamp 1018054153
transform 1 0 2896 0 1 1940
box -16 -6 32 210
use FILL  FILL_637
timestamp 1018054153
transform 1 0 2880 0 1 1940
box -16 -6 32 210
use FILL  FILL_638
timestamp 1018054153
transform 1 0 2368 0 1 1940
box -16 -6 32 210
use FILL  FILL_639
timestamp 1018054153
transform 1 0 1968 0 1 1940
box -16 -6 32 210
use FILL  FILL_640
timestamp 1018054153
transform 1 0 1952 0 1 1940
box -16 -6 32 210
use FILL  FILL_641
timestamp 1018054153
transform 1 0 1936 0 1 1940
box -16 -6 32 210
use FILL  FILL_642
timestamp 1018054153
transform 1 0 816 0 1 1940
box -16 -6 32 210
use FILL  FILL_643
timestamp 1018054153
transform 1 0 800 0 1 1940
box -16 -6 32 210
use FILL  FILL_644
timestamp 1018054153
transform 1 0 784 0 1 1940
box -16 -6 32 210
use FILL  FILL_645
timestamp 1018054153
transform 1 0 768 0 1 1940
box -16 -6 32 210
use FILL  FILL_646
timestamp 1018054153
transform 1 0 752 0 1 1940
box -16 -6 32 210
use FILL  FILL_647
timestamp 1018054153
transform 1 0 624 0 1 1940
box -16 -6 32 210
use FILL  FILL_648
timestamp 1018054153
transform 1 0 608 0 1 1940
box -16 -6 32 210
use FILL  FILL_649
timestamp 1018054153
transform 1 0 592 0 1 1940
box -16 -6 32 210
use FILL  FILL_650
timestamp 1018054153
transform 1 0 576 0 1 1940
box -16 -6 32 210
use FILL  FILL_651
timestamp 1018054153
transform 1 0 560 0 1 1940
box -16 -6 32 210
use FILL  FILL_652
timestamp 1018054153
transform 1 0 544 0 1 1940
box -16 -6 32 210
use FILL  FILL_653
timestamp 1018054153
transform 1 0 528 0 1 1940
box -16 -6 32 210
use FILL  FILL_654
timestamp 1018054153
transform 1 0 512 0 1 1940
box -16 -6 32 210
use FILL  FILL_655
timestamp 1018054153
transform 1 0 496 0 1 1940
box -16 -6 32 210
use FILL  FILL_656
timestamp 1018054153
transform 1 0 480 0 1 1940
box -16 -6 32 210
use FILL  FILL_657
timestamp 1018054153
transform 1 0 464 0 1 1940
box -16 -6 32 210
use FILL  FILL_658
timestamp 1018054153
transform 1 0 448 0 1 1940
box -16 -6 32 210
use FILL  FILL_659
timestamp 1018054153
transform 1 0 432 0 1 1940
box -16 -6 32 210
use FILL  FILL_660
timestamp 1018054153
transform 1 0 416 0 1 1940
box -16 -6 32 210
use FILL  FILL_661
timestamp 1018054153
transform 1 0 400 0 1 1940
box -16 -6 32 210
use FILL  FILL_662
timestamp 1018054153
transform 1 0 384 0 1 1940
box -16 -6 32 210
use FILL  FILL_663
timestamp 1018054153
transform 1 0 368 0 1 1940
box -16 -6 32 210
use FILL  FILL_664
timestamp 1018054153
transform 1 0 352 0 1 1940
box -16 -6 32 210
use FILL  FILL_665
timestamp 1018054153
transform 1 0 336 0 1 1940
box -16 -6 32 210
use FILL  FILL_666
timestamp 1018054153
transform 1 0 320 0 1 1940
box -16 -6 32 210
use FILL  FILL_667
timestamp 1018054153
transform 1 0 304 0 1 1940
box -16 -6 32 210
use FILL  FILL_668
timestamp 1018054153
transform 1 0 288 0 1 1940
box -16 -6 32 210
use FILL  FILL_669
timestamp 1018054153
transform 1 0 272 0 1 1940
box -16 -6 32 210
use FILL  FILL_670
timestamp 1018054153
transform 1 0 256 0 1 1940
box -16 -6 32 210
use FILL  FILL_671
timestamp 1018054153
transform 1 0 240 0 1 1940
box -16 -6 32 210
use FILL  FILL_672
timestamp 1018054153
transform 1 0 224 0 1 1940
box -16 -6 32 210
use FILL  FILL_673
timestamp 1018054153
transform 1 0 208 0 1 1940
box -16 -6 32 210
use FILL  FILL_674
timestamp 1018054153
transform 1 0 192 0 1 1940
box -16 -6 32 210
use FILL  FILL_675
timestamp 1018054153
transform 1 0 176 0 1 1940
box -16 -6 32 210
use FILL  FILL_676
timestamp 1018054153
transform 1 0 160 0 1 1940
box -16 -6 32 210
use FILL  FILL_677
timestamp 1018054153
transform 1 0 144 0 1 1940
box -16 -6 32 210
use FILL  FILL_678
timestamp 1018054153
transform 1 0 3664 0 -1 1940
box -16 -6 32 210
use FILL  FILL_679
timestamp 1018054153
transform 1 0 3648 0 -1 1940
box -16 -6 32 210
use FILL  FILL_680
timestamp 1018054153
transform 1 0 3632 0 -1 1940
box -16 -6 32 210
use FILL  FILL_681
timestamp 1018054153
transform 1 0 3616 0 -1 1940
box -16 -6 32 210
use FILL  FILL_682
timestamp 1018054153
transform 1 0 3600 0 -1 1940
box -16 -6 32 210
use FILL  FILL_683
timestamp 1018054153
transform 1 0 3584 0 -1 1940
box -16 -6 32 210
use FILL  FILL_684
timestamp 1018054153
transform 1 0 3568 0 -1 1940
box -16 -6 32 210
use FILL  FILL_685
timestamp 1018054153
transform 1 0 3552 0 -1 1940
box -16 -6 32 210
use FILL  FILL_686
timestamp 1018054153
transform 1 0 3536 0 -1 1940
box -16 -6 32 210
use FILL  FILL_687
timestamp 1018054153
transform 1 0 3520 0 -1 1940
box -16 -6 32 210
use FILL  FILL_688
timestamp 1018054153
transform 1 0 3504 0 -1 1940
box -16 -6 32 210
use FILL  FILL_689
timestamp 1018054153
transform 1 0 3200 0 -1 1940
box -16 -6 32 210
use FILL  FILL_690
timestamp 1018054153
transform 1 0 3184 0 -1 1940
box -16 -6 32 210
use FILL  FILL_691
timestamp 1018054153
transform 1 0 2976 0 -1 1940
box -16 -6 32 210
use FILL  FILL_692
timestamp 1018054153
transform 1 0 2960 0 -1 1940
box -16 -6 32 210
use FILL  FILL_693
timestamp 1018054153
transform 1 0 2944 0 -1 1940
box -16 -6 32 210
use FILL  FILL_694
timestamp 1018054153
transform 1 0 2928 0 -1 1940
box -16 -6 32 210
use FILL  FILL_695
timestamp 1018054153
transform 1 0 2912 0 -1 1940
box -16 -6 32 210
use FILL  FILL_696
timestamp 1018054153
transform 1 0 2800 0 -1 1940
box -16 -6 32 210
use FILL  FILL_697
timestamp 1018054153
transform 1 0 2784 0 -1 1940
box -16 -6 32 210
use FILL  FILL_698
timestamp 1018054153
transform 1 0 2576 0 -1 1940
box -16 -6 32 210
use FILL  FILL_699
timestamp 1018054153
transform 1 0 2560 0 -1 1940
box -16 -6 32 210
use FILL  FILL_700
timestamp 1018054153
transform 1 0 2544 0 -1 1940
box -16 -6 32 210
use FILL  FILL_701
timestamp 1018054153
transform 1 0 2528 0 -1 1940
box -16 -6 32 210
use FILL  FILL_702
timestamp 1018054153
transform 1 0 2400 0 -1 1940
box -16 -6 32 210
use FILL  FILL_703
timestamp 1018054153
transform 1 0 2384 0 -1 1940
box -16 -6 32 210
use FILL  FILL_704
timestamp 1018054153
transform 1 0 2368 0 -1 1940
box -16 -6 32 210
use FILL  FILL_705
timestamp 1018054153
transform 1 0 2352 0 -1 1940
box -16 -6 32 210
use FILL  FILL_706
timestamp 1018054153
transform 1 0 2336 0 -1 1940
box -16 -6 32 210
use FILL  FILL_707
timestamp 1018054153
transform 1 0 2320 0 -1 1940
box -16 -6 32 210
use FILL  FILL_708
timestamp 1018054153
transform 1 0 2208 0 -1 1940
box -16 -6 32 210
use FILL  FILL_709
timestamp 1018054153
transform 1 0 2192 0 -1 1940
box -16 -6 32 210
use FILL  FILL_710
timestamp 1018054153
transform 1 0 2176 0 -1 1940
box -16 -6 32 210
use FILL  FILL_711
timestamp 1018054153
transform 1 0 2160 0 -1 1940
box -16 -6 32 210
use FILL  FILL_712
timestamp 1018054153
transform 1 0 2144 0 -1 1940
box -16 -6 32 210
use FILL  FILL_713
timestamp 1018054153
transform 1 0 1904 0 -1 1940
box -16 -6 32 210
use FILL  FILL_714
timestamp 1018054153
transform 1 0 1888 0 -1 1940
box -16 -6 32 210
use FILL  FILL_715
timestamp 1018054153
transform 1 0 1872 0 -1 1940
box -16 -6 32 210
use FILL  FILL_716
timestamp 1018054153
transform 1 0 1856 0 -1 1940
box -16 -6 32 210
use FILL  FILL_717
timestamp 1018054153
transform 1 0 1840 0 -1 1940
box -16 -6 32 210
use FILL  FILL_718
timestamp 1018054153
transform 1 0 1824 0 -1 1940
box -16 -6 32 210
use FILL  FILL_719
timestamp 1018054153
transform 1 0 1808 0 -1 1940
box -16 -6 32 210
use FILL  FILL_720
timestamp 1018054153
transform 1 0 1792 0 -1 1940
box -16 -6 32 210
use FILL  FILL_721
timestamp 1018054153
transform 1 0 1664 0 -1 1940
box -16 -6 32 210
use FILL  FILL_722
timestamp 1018054153
transform 1 0 1648 0 -1 1940
box -16 -6 32 210
use FILL  FILL_723
timestamp 1018054153
transform 1 0 1632 0 -1 1940
box -16 -6 32 210
use FILL  FILL_724
timestamp 1018054153
transform 1 0 1424 0 -1 1940
box -16 -6 32 210
use FILL  FILL_725
timestamp 1018054153
transform 1 0 1408 0 -1 1940
box -16 -6 32 210
use FILL  FILL_726
timestamp 1018054153
transform 1 0 1392 0 -1 1940
box -16 -6 32 210
use FILL  FILL_727
timestamp 1018054153
transform 1 0 1376 0 -1 1940
box -16 -6 32 210
use FILL  FILL_728
timestamp 1018054153
transform 1 0 1360 0 -1 1940
box -16 -6 32 210
use FILL  FILL_729
timestamp 1018054153
transform 1 0 1264 0 -1 1940
box -16 -6 32 210
use FILL  FILL_730
timestamp 1018054153
transform 1 0 1248 0 -1 1940
box -16 -6 32 210
use FILL  FILL_731
timestamp 1018054153
transform 1 0 1232 0 -1 1940
box -16 -6 32 210
use FILL  FILL_732
timestamp 1018054153
transform 1 0 1024 0 -1 1940
box -16 -6 32 210
use FILL  FILL_733
timestamp 1018054153
transform 1 0 1008 0 -1 1940
box -16 -6 32 210
use FILL  FILL_734
timestamp 1018054153
transform 1 0 992 0 -1 1940
box -16 -6 32 210
use FILL  FILL_735
timestamp 1018054153
transform 1 0 912 0 -1 1940
box -16 -6 32 210
use FILL  FILL_736
timestamp 1018054153
transform 1 0 896 0 -1 1940
box -16 -6 32 210
use FILL  FILL_737
timestamp 1018054153
transform 1 0 880 0 -1 1940
box -16 -6 32 210
use FILL  FILL_738
timestamp 1018054153
transform 1 0 864 0 -1 1940
box -16 -6 32 210
use FILL  FILL_739
timestamp 1018054153
transform 1 0 848 0 -1 1940
box -16 -6 32 210
use FILL  FILL_740
timestamp 1018054153
transform 1 0 640 0 -1 1940
box -16 -6 32 210
use FILL  FILL_741
timestamp 1018054153
transform 1 0 576 0 -1 1940
box -16 -6 32 210
use FILL  FILL_742
timestamp 1018054153
transform 1 0 560 0 -1 1940
box -16 -6 32 210
use FILL  FILL_743
timestamp 1018054153
transform 1 0 544 0 -1 1940
box -16 -6 32 210
use FILL  FILL_744
timestamp 1018054153
transform 1 0 528 0 -1 1940
box -16 -6 32 210
use FILL  FILL_745
timestamp 1018054153
transform 1 0 512 0 -1 1940
box -16 -6 32 210
use FILL  FILL_746
timestamp 1018054153
transform 1 0 496 0 -1 1940
box -16 -6 32 210
use FILL  FILL_747
timestamp 1018054153
transform 1 0 480 0 -1 1940
box -16 -6 32 210
use FILL  FILL_748
timestamp 1018054153
transform 1 0 464 0 -1 1940
box -16 -6 32 210
use FILL  FILL_749
timestamp 1018054153
transform 1 0 448 0 -1 1940
box -16 -6 32 210
use FILL  FILL_750
timestamp 1018054153
transform 1 0 432 0 -1 1940
box -16 -6 32 210
use FILL  FILL_751
timestamp 1018054153
transform 1 0 416 0 -1 1940
box -16 -6 32 210
use FILL  FILL_752
timestamp 1018054153
transform 1 0 400 0 -1 1940
box -16 -6 32 210
use FILL  FILL_753
timestamp 1018054153
transform 1 0 384 0 -1 1940
box -16 -6 32 210
use FILL  FILL_754
timestamp 1018054153
transform 1 0 368 0 -1 1940
box -16 -6 32 210
use FILL  FILL_755
timestamp 1018054153
transform 1 0 352 0 -1 1940
box -16 -6 32 210
use FILL  FILL_756
timestamp 1018054153
transform 1 0 336 0 -1 1940
box -16 -6 32 210
use FILL  FILL_757
timestamp 1018054153
transform 1 0 320 0 -1 1940
box -16 -6 32 210
use FILL  FILL_758
timestamp 1018054153
transform 1 0 304 0 -1 1940
box -16 -6 32 210
use FILL  FILL_759
timestamp 1018054153
transform 1 0 288 0 -1 1940
box -16 -6 32 210
use FILL  FILL_760
timestamp 1018054153
transform 1 0 272 0 -1 1940
box -16 -6 32 210
use FILL  FILL_761
timestamp 1018054153
transform 1 0 256 0 -1 1940
box -16 -6 32 210
use FILL  FILL_762
timestamp 1018054153
transform 1 0 240 0 -1 1940
box -16 -6 32 210
use FILL  FILL_763
timestamp 1018054153
transform 1 0 224 0 -1 1940
box -16 -6 32 210
use FILL  FILL_764
timestamp 1018054153
transform 1 0 208 0 -1 1940
box -16 -6 32 210
use FILL  FILL_765
timestamp 1018054153
transform 1 0 192 0 -1 1940
box -16 -6 32 210
use FILL  FILL_766
timestamp 1018054153
transform 1 0 176 0 -1 1940
box -16 -6 32 210
use FILL  FILL_767
timestamp 1018054153
transform 1 0 160 0 -1 1940
box -16 -6 32 210
use FILL  FILL_768
timestamp 1018054153
transform 1 0 144 0 -1 1940
box -16 -6 32 210
use FILL  FILL_769
timestamp 1018054153
transform 1 0 3664 0 1 1540
box -16 -6 32 210
use FILL  FILL_770
timestamp 1018054153
transform 1 0 3648 0 1 1540
box -16 -6 32 210
use FILL  FILL_771
timestamp 1018054153
transform 1 0 3632 0 1 1540
box -16 -6 32 210
use FILL  FILL_772
timestamp 1018054153
transform 1 0 3616 0 1 1540
box -16 -6 32 210
use FILL  FILL_773
timestamp 1018054153
transform 1 0 3600 0 1 1540
box -16 -6 32 210
use FILL  FILL_774
timestamp 1018054153
transform 1 0 3584 0 1 1540
box -16 -6 32 210
use FILL  FILL_775
timestamp 1018054153
transform 1 0 3568 0 1 1540
box -16 -6 32 210
use FILL  FILL_776
timestamp 1018054153
transform 1 0 3552 0 1 1540
box -16 -6 32 210
use FILL  FILL_777
timestamp 1018054153
transform 1 0 3536 0 1 1540
box -16 -6 32 210
use FILL  FILL_778
timestamp 1018054153
transform 1 0 3520 0 1 1540
box -16 -6 32 210
use FILL  FILL_779
timestamp 1018054153
transform 1 0 3504 0 1 1540
box -16 -6 32 210
use FILL  FILL_780
timestamp 1018054153
transform 1 0 3280 0 1 1540
box -16 -6 32 210
use FILL  FILL_781
timestamp 1018054153
transform 1 0 3216 0 1 1540
box -16 -6 32 210
use FILL  FILL_782
timestamp 1018054153
transform 1 0 3200 0 1 1540
box -16 -6 32 210
use FILL  FILL_783
timestamp 1018054153
transform 1 0 3184 0 1 1540
box -16 -6 32 210
use FILL  FILL_784
timestamp 1018054153
transform 1 0 3168 0 1 1540
box -16 -6 32 210
use FILL  FILL_785
timestamp 1018054153
transform 1 0 3152 0 1 1540
box -16 -6 32 210
use FILL  FILL_786
timestamp 1018054153
transform 1 0 2816 0 1 1540
box -16 -6 32 210
use FILL  FILL_787
timestamp 1018054153
transform 1 0 2800 0 1 1540
box -16 -6 32 210
use FILL  FILL_788
timestamp 1018054153
transform 1 0 2784 0 1 1540
box -16 -6 32 210
use FILL  FILL_789
timestamp 1018054153
transform 1 0 2544 0 1 1540
box -16 -6 32 210
use FILL  FILL_790
timestamp 1018054153
transform 1 0 2416 0 1 1540
box -16 -6 32 210
use FILL  FILL_791
timestamp 1018054153
transform 1 0 2400 0 1 1540
box -16 -6 32 210
use FILL  FILL_792
timestamp 1018054153
transform 1 0 2384 0 1 1540
box -16 -6 32 210
use FILL  FILL_793
timestamp 1018054153
transform 1 0 2368 0 1 1540
box -16 -6 32 210
use FILL  FILL_794
timestamp 1018054153
transform 1 0 2352 0 1 1540
box -16 -6 32 210
use FILL  FILL_795
timestamp 1018054153
transform 1 0 2336 0 1 1540
box -16 -6 32 210
use FILL  FILL_796
timestamp 1018054153
transform 1 0 2320 0 1 1540
box -16 -6 32 210
use FILL  FILL_797
timestamp 1018054153
transform 1 0 2192 0 1 1540
box -16 -6 32 210
use FILL  FILL_798
timestamp 1018054153
transform 1 0 2176 0 1 1540
box -16 -6 32 210
use FILL  FILL_799
timestamp 1018054153
transform 1 0 2160 0 1 1540
box -16 -6 32 210
use FILL  FILL_800
timestamp 1018054153
transform 1 0 2144 0 1 1540
box -16 -6 32 210
use FILL  FILL_801
timestamp 1018054153
transform 1 0 2128 0 1 1540
box -16 -6 32 210
use FILL  FILL_802
timestamp 1018054153
transform 1 0 1664 0 1 1540
box -16 -6 32 210
use FILL  FILL_803
timestamp 1018054153
transform 1 0 1648 0 1 1540
box -16 -6 32 210
use FILL  FILL_804
timestamp 1018054153
transform 1 0 1632 0 1 1540
box -16 -6 32 210
use FILL  FILL_805
timestamp 1018054153
transform 1 0 1616 0 1 1540
box -16 -6 32 210
use FILL  FILL_806
timestamp 1018054153
transform 1 0 1600 0 1 1540
box -16 -6 32 210
use FILL  FILL_807
timestamp 1018054153
transform 1 0 1584 0 1 1540
box -16 -6 32 210
use FILL  FILL_808
timestamp 1018054153
transform 1 0 1264 0 1 1540
box -16 -6 32 210
use FILL  FILL_809
timestamp 1018054153
transform 1 0 1136 0 1 1540
box -16 -6 32 210
use FILL  FILL_810
timestamp 1018054153
transform 1 0 1120 0 1 1540
box -16 -6 32 210
use FILL  FILL_811
timestamp 1018054153
transform 1 0 1104 0 1 1540
box -16 -6 32 210
use FILL  FILL_812
timestamp 1018054153
transform 1 0 1088 0 1 1540
box -16 -6 32 210
use FILL  FILL_813
timestamp 1018054153
transform 1 0 1072 0 1 1540
box -16 -6 32 210
use FILL  FILL_814
timestamp 1018054153
transform 1 0 1056 0 1 1540
box -16 -6 32 210
use FILL  FILL_815
timestamp 1018054153
transform 1 0 1040 0 1 1540
box -16 -6 32 210
use FILL  FILL_816
timestamp 1018054153
transform 1 0 1024 0 1 1540
box -16 -6 32 210
use FILL  FILL_817
timestamp 1018054153
transform 1 0 944 0 1 1540
box -16 -6 32 210
use FILL  FILL_818
timestamp 1018054153
transform 1 0 928 0 1 1540
box -16 -6 32 210
use FILL  FILL_819
timestamp 1018054153
transform 1 0 912 0 1 1540
box -16 -6 32 210
use FILL  FILL_820
timestamp 1018054153
transform 1 0 848 0 1 1540
box -16 -6 32 210
use FILL  FILL_821
timestamp 1018054153
transform 1 0 800 0 1 1540
box -16 -6 32 210
use FILL  FILL_822
timestamp 1018054153
transform 1 0 784 0 1 1540
box -16 -6 32 210
use FILL  FILL_823
timestamp 1018054153
transform 1 0 768 0 1 1540
box -16 -6 32 210
use FILL  FILL_824
timestamp 1018054153
transform 1 0 752 0 1 1540
box -16 -6 32 210
use FILL  FILL_825
timestamp 1018054153
transform 1 0 736 0 1 1540
box -16 -6 32 210
use FILL  FILL_826
timestamp 1018054153
transform 1 0 720 0 1 1540
box -16 -6 32 210
use FILL  FILL_827
timestamp 1018054153
transform 1 0 704 0 1 1540
box -16 -6 32 210
use FILL  FILL_828
timestamp 1018054153
transform 1 0 544 0 1 1540
box -16 -6 32 210
use FILL  FILL_829
timestamp 1018054153
transform 1 0 528 0 1 1540
box -16 -6 32 210
use FILL  FILL_830
timestamp 1018054153
transform 1 0 512 0 1 1540
box -16 -6 32 210
use FILL  FILL_831
timestamp 1018054153
transform 1 0 496 0 1 1540
box -16 -6 32 210
use FILL  FILL_832
timestamp 1018054153
transform 1 0 480 0 1 1540
box -16 -6 32 210
use FILL  FILL_833
timestamp 1018054153
transform 1 0 464 0 1 1540
box -16 -6 32 210
use FILL  FILL_834
timestamp 1018054153
transform 1 0 448 0 1 1540
box -16 -6 32 210
use FILL  FILL_835
timestamp 1018054153
transform 1 0 432 0 1 1540
box -16 -6 32 210
use FILL  FILL_836
timestamp 1018054153
transform 1 0 416 0 1 1540
box -16 -6 32 210
use FILL  FILL_837
timestamp 1018054153
transform 1 0 400 0 1 1540
box -16 -6 32 210
use FILL  FILL_838
timestamp 1018054153
transform 1 0 384 0 1 1540
box -16 -6 32 210
use FILL  FILL_839
timestamp 1018054153
transform 1 0 368 0 1 1540
box -16 -6 32 210
use FILL  FILL_840
timestamp 1018054153
transform 1 0 352 0 1 1540
box -16 -6 32 210
use FILL  FILL_841
timestamp 1018054153
transform 1 0 336 0 1 1540
box -16 -6 32 210
use FILL  FILL_842
timestamp 1018054153
transform 1 0 320 0 1 1540
box -16 -6 32 210
use FILL  FILL_843
timestamp 1018054153
transform 1 0 304 0 1 1540
box -16 -6 32 210
use FILL  FILL_844
timestamp 1018054153
transform 1 0 288 0 1 1540
box -16 -6 32 210
use FILL  FILL_845
timestamp 1018054153
transform 1 0 272 0 1 1540
box -16 -6 32 210
use FILL  FILL_846
timestamp 1018054153
transform 1 0 256 0 1 1540
box -16 -6 32 210
use FILL  FILL_847
timestamp 1018054153
transform 1 0 240 0 1 1540
box -16 -6 32 210
use FILL  FILL_848
timestamp 1018054153
transform 1 0 224 0 1 1540
box -16 -6 32 210
use FILL  FILL_849
timestamp 1018054153
transform 1 0 208 0 1 1540
box -16 -6 32 210
use FILL  FILL_850
timestamp 1018054153
transform 1 0 192 0 1 1540
box -16 -6 32 210
use FILL  FILL_851
timestamp 1018054153
transform 1 0 176 0 1 1540
box -16 -6 32 210
use FILL  FILL_852
timestamp 1018054153
transform 1 0 160 0 1 1540
box -16 -6 32 210
use FILL  FILL_853
timestamp 1018054153
transform 1 0 144 0 1 1540
box -16 -6 32 210
use FILL  FILL_854
timestamp 1018054153
transform 1 0 3664 0 -1 1540
box -16 -6 32 210
use FILL  FILL_855
timestamp 1018054153
transform 1 0 3648 0 -1 1540
box -16 -6 32 210
use FILL  FILL_856
timestamp 1018054153
transform 1 0 3632 0 -1 1540
box -16 -6 32 210
use FILL  FILL_857
timestamp 1018054153
transform 1 0 3616 0 -1 1540
box -16 -6 32 210
use FILL  FILL_858
timestamp 1018054153
transform 1 0 3600 0 -1 1540
box -16 -6 32 210
use FILL  FILL_859
timestamp 1018054153
transform 1 0 3584 0 -1 1540
box -16 -6 32 210
use FILL  FILL_860
timestamp 1018054153
transform 1 0 3568 0 -1 1540
box -16 -6 32 210
use FILL  FILL_861
timestamp 1018054153
transform 1 0 3552 0 -1 1540
box -16 -6 32 210
use FILL  FILL_862
timestamp 1018054153
transform 1 0 3536 0 -1 1540
box -16 -6 32 210
use FILL  FILL_863
timestamp 1018054153
transform 1 0 3520 0 -1 1540
box -16 -6 32 210
use FILL  FILL_864
timestamp 1018054153
transform 1 0 3472 0 -1 1540
box -16 -6 32 210
use FILL  FILL_865
timestamp 1018054153
transform 1 0 3456 0 -1 1540
box -16 -6 32 210
use FILL  FILL_866
timestamp 1018054153
transform 1 0 3440 0 -1 1540
box -16 -6 32 210
use FILL  FILL_867
timestamp 1018054153
transform 1 0 3424 0 -1 1540
box -16 -6 32 210
use FILL  FILL_868
timestamp 1018054153
transform 1 0 3408 0 -1 1540
box -16 -6 32 210
use FILL  FILL_869
timestamp 1018054153
transform 1 0 3392 0 -1 1540
box -16 -6 32 210
use FILL  FILL_870
timestamp 1018054153
transform 1 0 3248 0 -1 1540
box -16 -6 32 210
use FILL  FILL_871
timestamp 1018054153
transform 1 0 3232 0 -1 1540
box -16 -6 32 210
use FILL  FILL_872
timestamp 1018054153
transform 1 0 2912 0 -1 1540
box -16 -6 32 210
use FILL  FILL_873
timestamp 1018054153
transform 1 0 2896 0 -1 1540
box -16 -6 32 210
use FILL  FILL_874
timestamp 1018054153
transform 1 0 2880 0 -1 1540
box -16 -6 32 210
use FILL  FILL_875
timestamp 1018054153
transform 1 0 2864 0 -1 1540
box -16 -6 32 210
use FILL  FILL_876
timestamp 1018054153
transform 1 0 2848 0 -1 1540
box -16 -6 32 210
use FILL  FILL_877
timestamp 1018054153
transform 1 0 2832 0 -1 1540
box -16 -6 32 210
use FILL  FILL_878
timestamp 1018054153
transform 1 0 2816 0 -1 1540
box -16 -6 32 210
use FILL  FILL_879
timestamp 1018054153
transform 1 0 2800 0 -1 1540
box -16 -6 32 210
use FILL  FILL_880
timestamp 1018054153
transform 1 0 2784 0 -1 1540
box -16 -6 32 210
use FILL  FILL_881
timestamp 1018054153
transform 1 0 2768 0 -1 1540
box -16 -6 32 210
use FILL  FILL_882
timestamp 1018054153
transform 1 0 2752 0 -1 1540
box -16 -6 32 210
use FILL  FILL_883
timestamp 1018054153
transform 1 0 2736 0 -1 1540
box -16 -6 32 210
use FILL  FILL_884
timestamp 1018054153
transform 1 0 2720 0 -1 1540
box -16 -6 32 210
use FILL  FILL_885
timestamp 1018054153
transform 1 0 2704 0 -1 1540
box -16 -6 32 210
use FILL  FILL_886
timestamp 1018054153
transform 1 0 1952 0 -1 1540
box -16 -6 32 210
use FILL  FILL_887
timestamp 1018054153
transform 1 0 1936 0 -1 1540
box -16 -6 32 210
use FILL  FILL_888
timestamp 1018054153
transform 1 0 1920 0 -1 1540
box -16 -6 32 210
use FILL  FILL_889
timestamp 1018054153
transform 1 0 1728 0 -1 1540
box -16 -6 32 210
use FILL  FILL_890
timestamp 1018054153
transform 1 0 1712 0 -1 1540
box -16 -6 32 210
use FILL  FILL_891
timestamp 1018054153
transform 1 0 1584 0 -1 1540
box -16 -6 32 210
use FILL  FILL_892
timestamp 1018054153
transform 1 0 1296 0 -1 1540
box -16 -6 32 210
use FILL  FILL_893
timestamp 1018054153
transform 1 0 1216 0 -1 1540
box -16 -6 32 210
use FILL  FILL_894
timestamp 1018054153
transform 1 0 1200 0 -1 1540
box -16 -6 32 210
use FILL  FILL_895
timestamp 1018054153
transform 1 0 1184 0 -1 1540
box -16 -6 32 210
use FILL  FILL_896
timestamp 1018054153
transform 1 0 1168 0 -1 1540
box -16 -6 32 210
use FILL  FILL_897
timestamp 1018054153
transform 1 0 1152 0 -1 1540
box -16 -6 32 210
use FILL  FILL_898
timestamp 1018054153
transform 1 0 1136 0 -1 1540
box -16 -6 32 210
use FILL  FILL_899
timestamp 1018054153
transform 1 0 1120 0 -1 1540
box -16 -6 32 210
use FILL  FILL_900
timestamp 1018054153
transform 1 0 992 0 -1 1540
box -16 -6 32 210
use FILL  FILL_901
timestamp 1018054153
transform 1 0 976 0 -1 1540
box -16 -6 32 210
use FILL  FILL_902
timestamp 1018054153
transform 1 0 928 0 -1 1540
box -16 -6 32 210
use FILL  FILL_903
timestamp 1018054153
transform 1 0 912 0 -1 1540
box -16 -6 32 210
use FILL  FILL_904
timestamp 1018054153
transform 1 0 896 0 -1 1540
box -16 -6 32 210
use FILL  FILL_905
timestamp 1018054153
transform 1 0 880 0 -1 1540
box -16 -6 32 210
use FILL  FILL_906
timestamp 1018054153
transform 1 0 864 0 -1 1540
box -16 -6 32 210
use FILL  FILL_907
timestamp 1018054153
transform 1 0 848 0 -1 1540
box -16 -6 32 210
use FILL  FILL_908
timestamp 1018054153
transform 1 0 832 0 -1 1540
box -16 -6 32 210
use FILL  FILL_909
timestamp 1018054153
transform 1 0 720 0 -1 1540
box -16 -6 32 210
use FILL  FILL_910
timestamp 1018054153
transform 1 0 704 0 -1 1540
box -16 -6 32 210
use FILL  FILL_911
timestamp 1018054153
transform 1 0 688 0 -1 1540
box -16 -6 32 210
use FILL  FILL_912
timestamp 1018054153
transform 1 0 672 0 -1 1540
box -16 -6 32 210
use FILL  FILL_913
timestamp 1018054153
transform 1 0 656 0 -1 1540
box -16 -6 32 210
use FILL  FILL_914
timestamp 1018054153
transform 1 0 640 0 -1 1540
box -16 -6 32 210
use FILL  FILL_915
timestamp 1018054153
transform 1 0 576 0 -1 1540
box -16 -6 32 210
use FILL  FILL_916
timestamp 1018054153
transform 1 0 560 0 -1 1540
box -16 -6 32 210
use FILL  FILL_917
timestamp 1018054153
transform 1 0 544 0 -1 1540
box -16 -6 32 210
use FILL  FILL_918
timestamp 1018054153
transform 1 0 528 0 -1 1540
box -16 -6 32 210
use FILL  FILL_919
timestamp 1018054153
transform 1 0 512 0 -1 1540
box -16 -6 32 210
use FILL  FILL_920
timestamp 1018054153
transform 1 0 496 0 -1 1540
box -16 -6 32 210
use FILL  FILL_921
timestamp 1018054153
transform 1 0 480 0 -1 1540
box -16 -6 32 210
use FILL  FILL_922
timestamp 1018054153
transform 1 0 464 0 -1 1540
box -16 -6 32 210
use FILL  FILL_923
timestamp 1018054153
transform 1 0 448 0 -1 1540
box -16 -6 32 210
use FILL  FILL_924
timestamp 1018054153
transform 1 0 432 0 -1 1540
box -16 -6 32 210
use FILL  FILL_925
timestamp 1018054153
transform 1 0 416 0 -1 1540
box -16 -6 32 210
use FILL  FILL_926
timestamp 1018054153
transform 1 0 400 0 -1 1540
box -16 -6 32 210
use FILL  FILL_927
timestamp 1018054153
transform 1 0 384 0 -1 1540
box -16 -6 32 210
use FILL  FILL_928
timestamp 1018054153
transform 1 0 368 0 -1 1540
box -16 -6 32 210
use FILL  FILL_929
timestamp 1018054153
transform 1 0 352 0 -1 1540
box -16 -6 32 210
use FILL  FILL_930
timestamp 1018054153
transform 1 0 336 0 -1 1540
box -16 -6 32 210
use FILL  FILL_931
timestamp 1018054153
transform 1 0 320 0 -1 1540
box -16 -6 32 210
use FILL  FILL_932
timestamp 1018054153
transform 1 0 304 0 -1 1540
box -16 -6 32 210
use FILL  FILL_933
timestamp 1018054153
transform 1 0 288 0 -1 1540
box -16 -6 32 210
use FILL  FILL_934
timestamp 1018054153
transform 1 0 272 0 -1 1540
box -16 -6 32 210
use FILL  FILL_935
timestamp 1018054153
transform 1 0 256 0 -1 1540
box -16 -6 32 210
use FILL  FILL_936
timestamp 1018054153
transform 1 0 240 0 -1 1540
box -16 -6 32 210
use FILL  FILL_937
timestamp 1018054153
transform 1 0 224 0 -1 1540
box -16 -6 32 210
use FILL  FILL_938
timestamp 1018054153
transform 1 0 208 0 -1 1540
box -16 -6 32 210
use FILL  FILL_939
timestamp 1018054153
transform 1 0 192 0 -1 1540
box -16 -6 32 210
use FILL  FILL_940
timestamp 1018054153
transform 1 0 176 0 -1 1540
box -16 -6 32 210
use FILL  FILL_941
timestamp 1018054153
transform 1 0 160 0 -1 1540
box -16 -6 32 210
use FILL  FILL_942
timestamp 1018054153
transform 1 0 144 0 -1 1540
box -16 -6 32 210
use FILL  FILL_943
timestamp 1018054153
transform 1 0 3424 0 1 1140
box -16 -6 32 210
use FILL  FILL_944
timestamp 1018054153
transform 1 0 3344 0 1 1140
box -16 -6 32 210
use FILL  FILL_945
timestamp 1018054153
transform 1 0 3328 0 1 1140
box -16 -6 32 210
use FILL  FILL_946
timestamp 1018054153
transform 1 0 3216 0 1 1140
box -16 -6 32 210
use FILL  FILL_947
timestamp 1018054153
transform 1 0 3200 0 1 1140
box -16 -6 32 210
use FILL  FILL_948
timestamp 1018054153
transform 1 0 3184 0 1 1140
box -16 -6 32 210
use FILL  FILL_949
timestamp 1018054153
transform 1 0 3168 0 1 1140
box -16 -6 32 210
use FILL  FILL_950
timestamp 1018054153
transform 1 0 2816 0 1 1140
box -16 -6 32 210
use FILL  FILL_951
timestamp 1018054153
transform 1 0 2800 0 1 1140
box -16 -6 32 210
use FILL  FILL_952
timestamp 1018054153
transform 1 0 2784 0 1 1140
box -16 -6 32 210
use FILL  FILL_953
timestamp 1018054153
transform 1 0 2768 0 1 1140
box -16 -6 32 210
use FILL  FILL_954
timestamp 1018054153
transform 1 0 2752 0 1 1140
box -16 -6 32 210
use FILL  FILL_955
timestamp 1018054153
transform 1 0 2288 0 1 1140
box -16 -6 32 210
use FILL  FILL_956
timestamp 1018054153
transform 1 0 2192 0 1 1140
box -16 -6 32 210
use FILL  FILL_957
timestamp 1018054153
transform 1 0 2176 0 1 1140
box -16 -6 32 210
use FILL  FILL_958
timestamp 1018054153
transform 1 0 2160 0 1 1140
box -16 -6 32 210
use FILL  FILL_959
timestamp 1018054153
transform 1 0 2144 0 1 1140
box -16 -6 32 210
use FILL  FILL_960
timestamp 1018054153
transform 1 0 1968 0 1 1140
box -16 -6 32 210
use FILL  FILL_961
timestamp 1018054153
transform 1 0 1648 0 1 1140
box -16 -6 32 210
use FILL  FILL_962
timestamp 1018054153
transform 1 0 1632 0 1 1140
box -16 -6 32 210
use FILL  FILL_963
timestamp 1018054153
transform 1 0 1616 0 1 1140
box -16 -6 32 210
use FILL  FILL_964
timestamp 1018054153
transform 1 0 1600 0 1 1140
box -16 -6 32 210
use FILL  FILL_965
timestamp 1018054153
transform 1 0 1584 0 1 1140
box -16 -6 32 210
use FILL  FILL_966
timestamp 1018054153
transform 1 0 1408 0 1 1140
box -16 -6 32 210
use FILL  FILL_967
timestamp 1018054153
transform 1 0 1392 0 1 1140
box -16 -6 32 210
use FILL  FILL_968
timestamp 1018054153
transform 1 0 1376 0 1 1140
box -16 -6 32 210
use FILL  FILL_969
timestamp 1018054153
transform 1 0 1360 0 1 1140
box -16 -6 32 210
use FILL  FILL_970
timestamp 1018054153
transform 1 0 1344 0 1 1140
box -16 -6 32 210
use FILL  FILL_971
timestamp 1018054153
transform 1 0 1328 0 1 1140
box -16 -6 32 210
use FILL  FILL_972
timestamp 1018054153
transform 1 0 1312 0 1 1140
box -16 -6 32 210
use FILL  FILL_973
timestamp 1018054153
transform 1 0 1296 0 1 1140
box -16 -6 32 210
use FILL  FILL_974
timestamp 1018054153
transform 1 0 1216 0 1 1140
box -16 -6 32 210
use FILL  FILL_975
timestamp 1018054153
transform 1 0 1200 0 1 1140
box -16 -6 32 210
use FILL  FILL_976
timestamp 1018054153
transform 1 0 1184 0 1 1140
box -16 -6 32 210
use FILL  FILL_977
timestamp 1018054153
transform 1 0 1168 0 1 1140
box -16 -6 32 210
use FILL  FILL_978
timestamp 1018054153
transform 1 0 1152 0 1 1140
box -16 -6 32 210
use FILL  FILL_979
timestamp 1018054153
transform 1 0 1136 0 1 1140
box -16 -6 32 210
use FILL  FILL_980
timestamp 1018054153
transform 1 0 1120 0 1 1140
box -16 -6 32 210
use FILL  FILL_981
timestamp 1018054153
transform 1 0 1056 0 1 1140
box -16 -6 32 210
use FILL  FILL_982
timestamp 1018054153
transform 1 0 1040 0 1 1140
box -16 -6 32 210
use FILL  FILL_983
timestamp 1018054153
transform 1 0 1024 0 1 1140
box -16 -6 32 210
use FILL  FILL_984
timestamp 1018054153
transform 1 0 1008 0 1 1140
box -16 -6 32 210
use FILL  FILL_985
timestamp 1018054153
transform 1 0 992 0 1 1140
box -16 -6 32 210
use FILL  FILL_986
timestamp 1018054153
transform 1 0 912 0 1 1140
box -16 -6 32 210
use FILL  FILL_987
timestamp 1018054153
transform 1 0 896 0 1 1140
box -16 -6 32 210
use FILL  FILL_988
timestamp 1018054153
transform 1 0 880 0 1 1140
box -16 -6 32 210
use FILL  FILL_989
timestamp 1018054153
transform 1 0 800 0 1 1140
box -16 -6 32 210
use FILL  FILL_990
timestamp 1018054153
transform 1 0 784 0 1 1140
box -16 -6 32 210
use FILL  FILL_991
timestamp 1018054153
transform 1 0 768 0 1 1140
box -16 -6 32 210
use FILL  FILL_992
timestamp 1018054153
transform 1 0 752 0 1 1140
box -16 -6 32 210
use FILL  FILL_993
timestamp 1018054153
transform 1 0 736 0 1 1140
box -16 -6 32 210
use FILL  FILL_994
timestamp 1018054153
transform 1 0 656 0 1 1140
box -16 -6 32 210
use FILL  FILL_995
timestamp 1018054153
transform 1 0 576 0 1 1140
box -16 -6 32 210
use FILL  FILL_996
timestamp 1018054153
transform 1 0 560 0 1 1140
box -16 -6 32 210
use FILL  FILL_997
timestamp 1018054153
transform 1 0 544 0 1 1140
box -16 -6 32 210
use FILL  FILL_998
timestamp 1018054153
transform 1 0 496 0 1 1140
box -16 -6 32 210
use FILL  FILL_999
timestamp 1018054153
transform 1 0 480 0 1 1140
box -16 -6 32 210
use FILL  FILL_1000
timestamp 1018054153
transform 1 0 464 0 1 1140
box -16 -6 32 210
use FILL  FILL_1001
timestamp 1018054153
transform 1 0 448 0 1 1140
box -16 -6 32 210
use FILL  FILL_1002
timestamp 1018054153
transform 1 0 432 0 1 1140
box -16 -6 32 210
use FILL  FILL_1003
timestamp 1018054153
transform 1 0 416 0 1 1140
box -16 -6 32 210
use FILL  FILL_1004
timestamp 1018054153
transform 1 0 400 0 1 1140
box -16 -6 32 210
use FILL  FILL_1005
timestamp 1018054153
transform 1 0 384 0 1 1140
box -16 -6 32 210
use FILL  FILL_1006
timestamp 1018054153
transform 1 0 368 0 1 1140
box -16 -6 32 210
use FILL  FILL_1007
timestamp 1018054153
transform 1 0 352 0 1 1140
box -16 -6 32 210
use FILL  FILL_1008
timestamp 1018054153
transform 1 0 336 0 1 1140
box -16 -6 32 210
use FILL  FILL_1009
timestamp 1018054153
transform 1 0 320 0 1 1140
box -16 -6 32 210
use FILL  FILL_1010
timestamp 1018054153
transform 1 0 304 0 1 1140
box -16 -6 32 210
use FILL  FILL_1011
timestamp 1018054153
transform 1 0 288 0 1 1140
box -16 -6 32 210
use FILL  FILL_1012
timestamp 1018054153
transform 1 0 272 0 1 1140
box -16 -6 32 210
use FILL  FILL_1013
timestamp 1018054153
transform 1 0 256 0 1 1140
box -16 -6 32 210
use FILL  FILL_1014
timestamp 1018054153
transform 1 0 240 0 1 1140
box -16 -6 32 210
use FILL  FILL_1015
timestamp 1018054153
transform 1 0 224 0 1 1140
box -16 -6 32 210
use FILL  FILL_1016
timestamp 1018054153
transform 1 0 208 0 1 1140
box -16 -6 32 210
use FILL  FILL_1017
timestamp 1018054153
transform 1 0 192 0 1 1140
box -16 -6 32 210
use FILL  FILL_1018
timestamp 1018054153
transform 1 0 176 0 1 1140
box -16 -6 32 210
use FILL  FILL_1019
timestamp 1018054153
transform 1 0 160 0 1 1140
box -16 -6 32 210
use FILL  FILL_1020
timestamp 1018054153
transform 1 0 144 0 1 1140
box -16 -6 32 210
use FILL  FILL_1021
timestamp 1018054153
transform 1 0 3664 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1022
timestamp 1018054153
transform 1 0 3648 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1023
timestamp 1018054153
transform 1 0 3632 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1024
timestamp 1018054153
transform 1 0 3616 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1025
timestamp 1018054153
transform 1 0 3440 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1026
timestamp 1018054153
transform 1 0 3424 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1027
timestamp 1018054153
transform 1 0 3408 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1028
timestamp 1018054153
transform 1 0 3392 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1029
timestamp 1018054153
transform 1 0 3248 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1030
timestamp 1018054153
transform 1 0 3232 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1031
timestamp 1018054153
transform 1 0 3216 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1032
timestamp 1018054153
transform 1 0 3200 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1033
timestamp 1018054153
transform 1 0 2736 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1034
timestamp 1018054153
transform 1 0 2720 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1035
timestamp 1018054153
transform 1 0 2704 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1036
timestamp 1018054153
transform 1 0 2688 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1037
timestamp 1018054153
transform 1 0 2560 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1038
timestamp 1018054153
transform 1 0 2544 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1039
timestamp 1018054153
transform 1 0 2528 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1040
timestamp 1018054153
transform 1 0 2320 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1041
timestamp 1018054153
transform 1 0 2304 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1042
timestamp 1018054153
transform 1 0 2288 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1043
timestamp 1018054153
transform 1 0 2160 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1044
timestamp 1018054153
transform 1 0 2144 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1045
timestamp 1018054153
transform 1 0 1968 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1046
timestamp 1018054153
transform 1 0 1952 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1047
timestamp 1018054153
transform 1 0 1904 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1048
timestamp 1018054153
transform 1 0 1888 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1049
timestamp 1018054153
transform 1 0 1872 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1050
timestamp 1018054153
transform 1 0 1856 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1051
timestamp 1018054153
transform 1 0 1840 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1052
timestamp 1018054153
transform 1 0 1824 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1053
timestamp 1018054153
transform 1 0 1808 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1054
timestamp 1018054153
transform 1 0 1680 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1055
timestamp 1018054153
transform 1 0 1664 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1056
timestamp 1018054153
transform 1 0 1648 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1057
timestamp 1018054153
transform 1 0 1632 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1058
timestamp 1018054153
transform 1 0 1616 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1059
timestamp 1018054153
transform 1 0 1424 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1060
timestamp 1018054153
transform 1 0 1408 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1061
timestamp 1018054153
transform 1 0 1392 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1062
timestamp 1018054153
transform 1 0 1376 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1063
timestamp 1018054153
transform 1 0 1360 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1064
timestamp 1018054153
transform 1 0 1232 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1065
timestamp 1018054153
transform 1 0 1216 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1066
timestamp 1018054153
transform 1 0 1200 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1067
timestamp 1018054153
transform 1 0 1120 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1068
timestamp 1018054153
transform 1 0 1040 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1069
timestamp 1018054153
transform 1 0 1024 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1070
timestamp 1018054153
transform 1 0 1008 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1071
timestamp 1018054153
transform 1 0 944 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1072
timestamp 1018054153
transform 1 0 880 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1073
timestamp 1018054153
transform 1 0 864 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1074
timestamp 1018054153
transform 1 0 848 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1075
timestamp 1018054153
transform 1 0 832 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1076
timestamp 1018054153
transform 1 0 816 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1077
timestamp 1018054153
transform 1 0 800 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1078
timestamp 1018054153
transform 1 0 656 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1079
timestamp 1018054153
transform 1 0 640 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1080
timestamp 1018054153
transform 1 0 624 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1081
timestamp 1018054153
transform 1 0 608 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1082
timestamp 1018054153
transform 1 0 592 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1083
timestamp 1018054153
transform 1 0 576 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1084
timestamp 1018054153
transform 1 0 304 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1085
timestamp 1018054153
transform 1 0 288 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1086
timestamp 1018054153
transform 1 0 272 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1087
timestamp 1018054153
transform 1 0 256 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1088
timestamp 1018054153
transform 1 0 240 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1089
timestamp 1018054153
transform 1 0 224 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1090
timestamp 1018054153
transform 1 0 208 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1091
timestamp 1018054153
transform 1 0 192 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1092
timestamp 1018054153
transform 1 0 176 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1093
timestamp 1018054153
transform 1 0 160 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1094
timestamp 1018054153
transform 1 0 144 0 -1 1140
box -16 -6 32 210
use FILL  FILL_1095
timestamp 1018054153
transform 1 0 3664 0 1 740
box -16 -6 32 210
use FILL  FILL_1096
timestamp 1018054153
transform 1 0 3648 0 1 740
box -16 -6 32 210
use FILL  FILL_1097
timestamp 1018054153
transform 1 0 3632 0 1 740
box -16 -6 32 210
use FILL  FILL_1098
timestamp 1018054153
transform 1 0 3616 0 1 740
box -16 -6 32 210
use FILL  FILL_1099
timestamp 1018054153
transform 1 0 3600 0 1 740
box -16 -6 32 210
use FILL  FILL_1100
timestamp 1018054153
transform 1 0 3584 0 1 740
box -16 -6 32 210
use FILL  FILL_1101
timestamp 1018054153
transform 1 0 3472 0 1 740
box -16 -6 32 210
use FILL  FILL_1102
timestamp 1018054153
transform 1 0 3456 0 1 740
box -16 -6 32 210
use FILL  FILL_1103
timestamp 1018054153
transform 1 0 3440 0 1 740
box -16 -6 32 210
use FILL  FILL_1104
timestamp 1018054153
transform 1 0 3424 0 1 740
box -16 -6 32 210
use FILL  FILL_1105
timestamp 1018054153
transform 1 0 3408 0 1 740
box -16 -6 32 210
use FILL  FILL_1106
timestamp 1018054153
transform 1 0 3392 0 1 740
box -16 -6 32 210
use FILL  FILL_1107
timestamp 1018054153
transform 1 0 3248 0 1 740
box -16 -6 32 210
use FILL  FILL_1108
timestamp 1018054153
transform 1 0 3232 0 1 740
box -16 -6 32 210
use FILL  FILL_1109
timestamp 1018054153
transform 1 0 3216 0 1 740
box -16 -6 32 210
use FILL  FILL_1110
timestamp 1018054153
transform 1 0 2560 0 1 740
box -16 -6 32 210
use FILL  FILL_1111
timestamp 1018054153
transform 1 0 2544 0 1 740
box -16 -6 32 210
use FILL  FILL_1112
timestamp 1018054153
transform 1 0 2528 0 1 740
box -16 -6 32 210
use FILL  FILL_1113
timestamp 1018054153
transform 1 0 2512 0 1 740
box -16 -6 32 210
use FILL  FILL_1114
timestamp 1018054153
transform 1 0 2416 0 1 740
box -16 -6 32 210
use FILL  FILL_1115
timestamp 1018054153
transform 1 0 2400 0 1 740
box -16 -6 32 210
use FILL  FILL_1116
timestamp 1018054153
transform 1 0 2384 0 1 740
box -16 -6 32 210
use FILL  FILL_1117
timestamp 1018054153
transform 1 0 2144 0 1 740
box -16 -6 32 210
use FILL  FILL_1118
timestamp 1018054153
transform 1 0 2128 0 1 740
box -16 -6 32 210
use FILL  FILL_1119
timestamp 1018054153
transform 1 0 2112 0 1 740
box -16 -6 32 210
use FILL  FILL_1120
timestamp 1018054153
transform 1 0 1856 0 1 740
box -16 -6 32 210
use FILL  FILL_1121
timestamp 1018054153
transform 1 0 1648 0 1 740
box -16 -6 32 210
use FILL  FILL_1122
timestamp 1018054153
transform 1 0 1632 0 1 740
box -16 -6 32 210
use FILL  FILL_1123
timestamp 1018054153
transform 1 0 1616 0 1 740
box -16 -6 32 210
use FILL  FILL_1124
timestamp 1018054153
transform 1 0 1552 0 1 740
box -16 -6 32 210
use FILL  FILL_1125
timestamp 1018054153
transform 1 0 1536 0 1 740
box -16 -6 32 210
use FILL  FILL_1126
timestamp 1018054153
transform 1 0 1520 0 1 740
box -16 -6 32 210
use FILL  FILL_1127
timestamp 1018054153
transform 1 0 1504 0 1 740
box -16 -6 32 210
use FILL  FILL_1128
timestamp 1018054153
transform 1 0 1488 0 1 740
box -16 -6 32 210
use FILL  FILL_1129
timestamp 1018054153
transform 1 0 1472 0 1 740
box -16 -6 32 210
use FILL  FILL_1130
timestamp 1018054153
transform 1 0 1456 0 1 740
box -16 -6 32 210
use FILL  FILL_1131
timestamp 1018054153
transform 1 0 1376 0 1 740
box -16 -6 32 210
use FILL  FILL_1132
timestamp 1018054153
transform 1 0 1360 0 1 740
box -16 -6 32 210
use FILL  FILL_1133
timestamp 1018054153
transform 1 0 1344 0 1 740
box -16 -6 32 210
use FILL  FILL_1134
timestamp 1018054153
transform 1 0 1328 0 1 740
box -16 -6 32 210
use FILL  FILL_1135
timestamp 1018054153
transform 1 0 1280 0 1 740
box -16 -6 32 210
use FILL  FILL_1136
timestamp 1018054153
transform 1 0 1232 0 1 740
box -16 -6 32 210
use FILL  FILL_1137
timestamp 1018054153
transform 1 0 1216 0 1 740
box -16 -6 32 210
use FILL  FILL_1138
timestamp 1018054153
transform 1 0 1200 0 1 740
box -16 -6 32 210
use FILL  FILL_1139
timestamp 1018054153
transform 1 0 1184 0 1 740
box -16 -6 32 210
use FILL  FILL_1140
timestamp 1018054153
transform 1 0 1168 0 1 740
box -16 -6 32 210
use FILL  FILL_1141
timestamp 1018054153
transform 1 0 1152 0 1 740
box -16 -6 32 210
use FILL  FILL_1142
timestamp 1018054153
transform 1 0 1136 0 1 740
box -16 -6 32 210
use FILL  FILL_1143
timestamp 1018054153
transform 1 0 1056 0 1 740
box -16 -6 32 210
use FILL  FILL_1144
timestamp 1018054153
transform 1 0 1040 0 1 740
box -16 -6 32 210
use FILL  FILL_1145
timestamp 1018054153
transform 1 0 1024 0 1 740
box -16 -6 32 210
use FILL  FILL_1146
timestamp 1018054153
transform 1 0 1008 0 1 740
box -16 -6 32 210
use FILL  FILL_1147
timestamp 1018054153
transform 1 0 992 0 1 740
box -16 -6 32 210
use FILL  FILL_1148
timestamp 1018054153
transform 1 0 880 0 1 740
box -16 -6 32 210
use FILL  FILL_1149
timestamp 1018054153
transform 1 0 864 0 1 740
box -16 -6 32 210
use FILL  FILL_1150
timestamp 1018054153
transform 1 0 848 0 1 740
box -16 -6 32 210
use FILL  FILL_1151
timestamp 1018054153
transform 1 0 832 0 1 740
box -16 -6 32 210
use FILL  FILL_1152
timestamp 1018054153
transform 1 0 816 0 1 740
box -16 -6 32 210
use FILL  FILL_1153
timestamp 1018054153
transform 1 0 800 0 1 740
box -16 -6 32 210
use FILL  FILL_1154
timestamp 1018054153
transform 1 0 688 0 1 740
box -16 -6 32 210
use FILL  FILL_1155
timestamp 1018054153
transform 1 0 672 0 1 740
box -16 -6 32 210
use FILL  FILL_1156
timestamp 1018054153
transform 1 0 608 0 1 740
box -16 -6 32 210
use FILL  FILL_1157
timestamp 1018054153
transform 1 0 592 0 1 740
box -16 -6 32 210
use FILL  FILL_1158
timestamp 1018054153
transform 1 0 576 0 1 740
box -16 -6 32 210
use FILL  FILL_1159
timestamp 1018054153
transform 1 0 560 0 1 740
box -16 -6 32 210
use FILL  FILL_1160
timestamp 1018054153
transform 1 0 432 0 1 740
box -16 -6 32 210
use FILL  FILL_1161
timestamp 1018054153
transform 1 0 416 0 1 740
box -16 -6 32 210
use FILL  FILL_1162
timestamp 1018054153
transform 1 0 400 0 1 740
box -16 -6 32 210
use FILL  FILL_1163
timestamp 1018054153
transform 1 0 384 0 1 740
box -16 -6 32 210
use FILL  FILL_1164
timestamp 1018054153
transform 1 0 368 0 1 740
box -16 -6 32 210
use FILL  FILL_1165
timestamp 1018054153
transform 1 0 352 0 1 740
box -16 -6 32 210
use FILL  FILL_1166
timestamp 1018054153
transform 1 0 336 0 1 740
box -16 -6 32 210
use FILL  FILL_1167
timestamp 1018054153
transform 1 0 320 0 1 740
box -16 -6 32 210
use FILL  FILL_1168
timestamp 1018054153
transform 1 0 304 0 1 740
box -16 -6 32 210
use FILL  FILL_1169
timestamp 1018054153
transform 1 0 288 0 1 740
box -16 -6 32 210
use FILL  FILL_1170
timestamp 1018054153
transform 1 0 272 0 1 740
box -16 -6 32 210
use FILL  FILL_1171
timestamp 1018054153
transform 1 0 256 0 1 740
box -16 -6 32 210
use FILL  FILL_1172
timestamp 1018054153
transform 1 0 240 0 1 740
box -16 -6 32 210
use FILL  FILL_1173
timestamp 1018054153
transform 1 0 224 0 1 740
box -16 -6 32 210
use FILL  FILL_1174
timestamp 1018054153
transform 1 0 208 0 1 740
box -16 -6 32 210
use FILL  FILL_1175
timestamp 1018054153
transform 1 0 192 0 1 740
box -16 -6 32 210
use FILL  FILL_1176
timestamp 1018054153
transform 1 0 176 0 1 740
box -16 -6 32 210
use FILL  FILL_1177
timestamp 1018054153
transform 1 0 160 0 1 740
box -16 -6 32 210
use FILL  FILL_1178
timestamp 1018054153
transform 1 0 144 0 1 740
box -16 -6 32 210
use FILL  FILL_1179
timestamp 1018054153
transform 1 0 3664 0 -1 740
box -16 -6 32 210
use FILL  FILL_1180
timestamp 1018054153
transform 1 0 3648 0 -1 740
box -16 -6 32 210
use FILL  FILL_1181
timestamp 1018054153
transform 1 0 3632 0 -1 740
box -16 -6 32 210
use FILL  FILL_1182
timestamp 1018054153
transform 1 0 3616 0 -1 740
box -16 -6 32 210
use FILL  FILL_1183
timestamp 1018054153
transform 1 0 3600 0 -1 740
box -16 -6 32 210
use FILL  FILL_1184
timestamp 1018054153
transform 1 0 3232 0 -1 740
box -16 -6 32 210
use FILL  FILL_1185
timestamp 1018054153
transform 1 0 2928 0 -1 740
box -16 -6 32 210
use FILL  FILL_1186
timestamp 1018054153
transform 1 0 2752 0 -1 740
box -16 -6 32 210
use FILL  FILL_1187
timestamp 1018054153
transform 1 0 2496 0 -1 740
box -16 -6 32 210
use FILL  FILL_1188
timestamp 1018054153
transform 1 0 2480 0 -1 740
box -16 -6 32 210
use FILL  FILL_1189
timestamp 1018054153
transform 1 0 2464 0 -1 740
box -16 -6 32 210
use FILL  FILL_1190
timestamp 1018054153
transform 1 0 2448 0 -1 740
box -16 -6 32 210
use FILL  FILL_1191
timestamp 1018054153
transform 1 0 2304 0 -1 740
box -16 -6 32 210
use FILL  FILL_1192
timestamp 1018054153
transform 1 0 2288 0 -1 740
box -16 -6 32 210
use FILL  FILL_1193
timestamp 1018054153
transform 1 0 2272 0 -1 740
box -16 -6 32 210
use FILL  FILL_1194
timestamp 1018054153
transform 1 0 2256 0 -1 740
box -16 -6 32 210
use FILL  FILL_1195
timestamp 1018054153
transform 1 0 2208 0 -1 740
box -16 -6 32 210
use FILL  FILL_1196
timestamp 1018054153
transform 1 0 2192 0 -1 740
box -16 -6 32 210
use FILL  FILL_1197
timestamp 1018054153
transform 1 0 2176 0 -1 740
box -16 -6 32 210
use FILL  FILL_1198
timestamp 1018054153
transform 1 0 2160 0 -1 740
box -16 -6 32 210
use FILL  FILL_1199
timestamp 1018054153
transform 1 0 2032 0 -1 740
box -16 -6 32 210
use FILL  FILL_1200
timestamp 1018054153
transform 1 0 2016 0 -1 740
box -16 -6 32 210
use FILL  FILL_1201
timestamp 1018054153
transform 1 0 2000 0 -1 740
box -16 -6 32 210
use FILL  FILL_1202
timestamp 1018054153
transform 1 0 1984 0 -1 740
box -16 -6 32 210
use FILL  FILL_1203
timestamp 1018054153
transform 1 0 1968 0 -1 740
box -16 -6 32 210
use FILL  FILL_1204
timestamp 1018054153
transform 1 0 1872 0 -1 740
box -16 -6 32 210
use FILL  FILL_1205
timestamp 1018054153
transform 1 0 1856 0 -1 740
box -16 -6 32 210
use FILL  FILL_1206
timestamp 1018054153
transform 1 0 1840 0 -1 740
box -16 -6 32 210
use FILL  FILL_1207
timestamp 1018054153
transform 1 0 1824 0 -1 740
box -16 -6 32 210
use FILL  FILL_1208
timestamp 1018054153
transform 1 0 1808 0 -1 740
box -16 -6 32 210
use FILL  FILL_1209
timestamp 1018054153
transform 1 0 1360 0 -1 740
box -16 -6 32 210
use FILL  FILL_1210
timestamp 1018054153
transform 1 0 1344 0 -1 740
box -16 -6 32 210
use FILL  FILL_1211
timestamp 1018054153
transform 1 0 1328 0 -1 740
box -16 -6 32 210
use FILL  FILL_1212
timestamp 1018054153
transform 1 0 1280 0 -1 740
box -16 -6 32 210
use FILL  FILL_1213
timestamp 1018054153
transform 1 0 1264 0 -1 740
box -16 -6 32 210
use FILL  FILL_1214
timestamp 1018054153
transform 1 0 1248 0 -1 740
box -16 -6 32 210
use FILL  FILL_1215
timestamp 1018054153
transform 1 0 1232 0 -1 740
box -16 -6 32 210
use FILL  FILL_1216
timestamp 1018054153
transform 1 0 1088 0 -1 740
box -16 -6 32 210
use FILL  FILL_1217
timestamp 1018054153
transform 1 0 1072 0 -1 740
box -16 -6 32 210
use FILL  FILL_1218
timestamp 1018054153
transform 1 0 1056 0 -1 740
box -16 -6 32 210
use FILL  FILL_1219
timestamp 1018054153
transform 1 0 1040 0 -1 740
box -16 -6 32 210
use FILL  FILL_1220
timestamp 1018054153
transform 1 0 1024 0 -1 740
box -16 -6 32 210
use FILL  FILL_1221
timestamp 1018054153
transform 1 0 1008 0 -1 740
box -16 -6 32 210
use FILL  FILL_1222
timestamp 1018054153
transform 1 0 992 0 -1 740
box -16 -6 32 210
use FILL  FILL_1223
timestamp 1018054153
transform 1 0 864 0 -1 740
box -16 -6 32 210
use FILL  FILL_1224
timestamp 1018054153
transform 1 0 848 0 -1 740
box -16 -6 32 210
use FILL  FILL_1225
timestamp 1018054153
transform 1 0 832 0 -1 740
box -16 -6 32 210
use FILL  FILL_1226
timestamp 1018054153
transform 1 0 816 0 -1 740
box -16 -6 32 210
use FILL  FILL_1227
timestamp 1018054153
transform 1 0 800 0 -1 740
box -16 -6 32 210
use FILL  FILL_1228
timestamp 1018054153
transform 1 0 784 0 -1 740
box -16 -6 32 210
use FILL  FILL_1229
timestamp 1018054153
transform 1 0 768 0 -1 740
box -16 -6 32 210
use FILL  FILL_1230
timestamp 1018054153
transform 1 0 656 0 -1 740
box -16 -6 32 210
use FILL  FILL_1231
timestamp 1018054153
transform 1 0 640 0 -1 740
box -16 -6 32 210
use FILL  FILL_1232
timestamp 1018054153
transform 1 0 624 0 -1 740
box -16 -6 32 210
use FILL  FILL_1233
timestamp 1018054153
transform 1 0 608 0 -1 740
box -16 -6 32 210
use FILL  FILL_1234
timestamp 1018054153
transform 1 0 592 0 -1 740
box -16 -6 32 210
use FILL  FILL_1235
timestamp 1018054153
transform 1 0 304 0 -1 740
box -16 -6 32 210
use FILL  FILL_1236
timestamp 1018054153
transform 1 0 288 0 -1 740
box -16 -6 32 210
use FILL  FILL_1237
timestamp 1018054153
transform 1 0 272 0 -1 740
box -16 -6 32 210
use FILL  FILL_1238
timestamp 1018054153
transform 1 0 256 0 -1 740
box -16 -6 32 210
use FILL  FILL_1239
timestamp 1018054153
transform 1 0 240 0 -1 740
box -16 -6 32 210
use FILL  FILL_1240
timestamp 1018054153
transform 1 0 224 0 -1 740
box -16 -6 32 210
use FILL  FILL_1241
timestamp 1018054153
transform 1 0 208 0 -1 740
box -16 -6 32 210
use FILL  FILL_1242
timestamp 1018054153
transform 1 0 192 0 -1 740
box -16 -6 32 210
use FILL  FILL_1243
timestamp 1018054153
transform 1 0 176 0 -1 740
box -16 -6 32 210
use FILL  FILL_1244
timestamp 1018054153
transform 1 0 160 0 -1 740
box -16 -6 32 210
use FILL  FILL_1245
timestamp 1018054153
transform 1 0 144 0 -1 740
box -16 -6 32 210
use FILL  FILL_1246
timestamp 1018054153
transform 1 0 3664 0 1 340
box -16 -6 32 210
use FILL  FILL_1247
timestamp 1018054153
transform 1 0 3648 0 1 340
box -16 -6 32 210
use FILL  FILL_1248
timestamp 1018054153
transform 1 0 3632 0 1 340
box -16 -6 32 210
use FILL  FILL_1249
timestamp 1018054153
transform 1 0 3408 0 1 340
box -16 -6 32 210
use FILL  FILL_1250
timestamp 1018054153
transform 1 0 3392 0 1 340
box -16 -6 32 210
use FILL  FILL_1251
timestamp 1018054153
transform 1 0 3376 0 1 340
box -16 -6 32 210
use FILL  FILL_1252
timestamp 1018054153
transform 1 0 3232 0 1 340
box -16 -6 32 210
use FILL  FILL_1253
timestamp 1018054153
transform 1 0 3216 0 1 340
box -16 -6 32 210
use FILL  FILL_1254
timestamp 1018054153
transform 1 0 3200 0 1 340
box -16 -6 32 210
use FILL  FILL_1255
timestamp 1018054153
transform 1 0 3184 0 1 340
box -16 -6 32 210
use FILL  FILL_1256
timestamp 1018054153
transform 1 0 3168 0 1 340
box -16 -6 32 210
use FILL  FILL_1257
timestamp 1018054153
transform 1 0 3056 0 1 340
box -16 -6 32 210
use FILL  FILL_1258
timestamp 1018054153
transform 1 0 3040 0 1 340
box -16 -6 32 210
use FILL  FILL_1259
timestamp 1018054153
transform 1 0 3024 0 1 340
box -16 -6 32 210
use FILL  FILL_1260
timestamp 1018054153
transform 1 0 2800 0 1 340
box -16 -6 32 210
use FILL  FILL_1261
timestamp 1018054153
transform 1 0 2784 0 1 340
box -16 -6 32 210
use FILL  FILL_1262
timestamp 1018054153
transform 1 0 2768 0 1 340
box -16 -6 32 210
use FILL  FILL_1263
timestamp 1018054153
transform 1 0 2752 0 1 340
box -16 -6 32 210
use FILL  FILL_1264
timestamp 1018054153
transform 1 0 2736 0 1 340
box -16 -6 32 210
use FILL  FILL_1265
timestamp 1018054153
transform 1 0 2720 0 1 340
box -16 -6 32 210
use FILL  FILL_1266
timestamp 1018054153
transform 1 0 2608 0 1 340
box -16 -6 32 210
use FILL  FILL_1267
timestamp 1018054153
transform 1 0 2592 0 1 340
box -16 -6 32 210
use FILL  FILL_1268
timestamp 1018054153
transform 1 0 2576 0 1 340
box -16 -6 32 210
use FILL  FILL_1269
timestamp 1018054153
transform 1 0 2560 0 1 340
box -16 -6 32 210
use FILL  FILL_1270
timestamp 1018054153
transform 1 0 2544 0 1 340
box -16 -6 32 210
use FILL  FILL_1271
timestamp 1018054153
transform 1 0 2480 0 1 340
box -16 -6 32 210
use FILL  FILL_1272
timestamp 1018054153
transform 1 0 2256 0 1 340
box -16 -6 32 210
use FILL  FILL_1273
timestamp 1018054153
transform 1 0 2240 0 1 340
box -16 -6 32 210
use FILL  FILL_1274
timestamp 1018054153
transform 1 0 2224 0 1 340
box -16 -6 32 210
use FILL  FILL_1275
timestamp 1018054153
transform 1 0 2208 0 1 340
box -16 -6 32 210
use FILL  FILL_1276
timestamp 1018054153
transform 1 0 2160 0 1 340
box -16 -6 32 210
use FILL  FILL_1277
timestamp 1018054153
transform 1 0 2144 0 1 340
box -16 -6 32 210
use FILL  FILL_1278
timestamp 1018054153
transform 1 0 2128 0 1 340
box -16 -6 32 210
use FILL  FILL_1279
timestamp 1018054153
transform 1 0 2112 0 1 340
box -16 -6 32 210
use FILL  FILL_1280
timestamp 1018054153
transform 1 0 2096 0 1 340
box -16 -6 32 210
use FILL  FILL_1281
timestamp 1018054153
transform 1 0 2080 0 1 340
box -16 -6 32 210
use FILL  FILL_1282
timestamp 1018054153
transform 1 0 2064 0 1 340
box -16 -6 32 210
use FILL  FILL_1283
timestamp 1018054153
transform 1 0 1600 0 1 340
box -16 -6 32 210
use FILL  FILL_1284
timestamp 1018054153
transform 1 0 1584 0 1 340
box -16 -6 32 210
use FILL  FILL_1285
timestamp 1018054153
transform 1 0 1568 0 1 340
box -16 -6 32 210
use FILL  FILL_1286
timestamp 1018054153
transform 1 0 1552 0 1 340
box -16 -6 32 210
use FILL  FILL_1287
timestamp 1018054153
transform 1 0 1536 0 1 340
box -16 -6 32 210
use FILL  FILL_1288
timestamp 1018054153
transform 1 0 1424 0 1 340
box -16 -6 32 210
use FILL  FILL_1289
timestamp 1018054153
transform 1 0 1408 0 1 340
box -16 -6 32 210
use FILL  FILL_1290
timestamp 1018054153
transform 1 0 1392 0 1 340
box -16 -6 32 210
use FILL  FILL_1291
timestamp 1018054153
transform 1 0 1376 0 1 340
box -16 -6 32 210
use FILL  FILL_1292
timestamp 1018054153
transform 1 0 1360 0 1 340
box -16 -6 32 210
use FILL  FILL_1293
timestamp 1018054153
transform 1 0 1344 0 1 340
box -16 -6 32 210
use FILL  FILL_1294
timestamp 1018054153
transform 1 0 1136 0 1 340
box -16 -6 32 210
use FILL  FILL_1295
timestamp 1018054153
transform 1 0 1120 0 1 340
box -16 -6 32 210
use FILL  FILL_1296
timestamp 1018054153
transform 1 0 1104 0 1 340
box -16 -6 32 210
use FILL  FILL_1297
timestamp 1018054153
transform 1 0 1088 0 1 340
box -16 -6 32 210
use FILL  FILL_1298
timestamp 1018054153
transform 1 0 1072 0 1 340
box -16 -6 32 210
use FILL  FILL_1299
timestamp 1018054153
transform 1 0 1056 0 1 340
box -16 -6 32 210
use FILL  FILL_1300
timestamp 1018054153
transform 1 0 1040 0 1 340
box -16 -6 32 210
use FILL  FILL_1301
timestamp 1018054153
transform 1 0 1024 0 1 340
box -16 -6 32 210
use FILL  FILL_1302
timestamp 1018054153
transform 1 0 1008 0 1 340
box -16 -6 32 210
use FILL  FILL_1303
timestamp 1018054153
transform 1 0 992 0 1 340
box -16 -6 32 210
use FILL  FILL_1304
timestamp 1018054153
transform 1 0 976 0 1 340
box -16 -6 32 210
use FILL  FILL_1305
timestamp 1018054153
transform 1 0 960 0 1 340
box -16 -6 32 210
use FILL  FILL_1306
timestamp 1018054153
transform 1 0 944 0 1 340
box -16 -6 32 210
use FILL  FILL_1307
timestamp 1018054153
transform 1 0 928 0 1 340
box -16 -6 32 210
use FILL  FILL_1308
timestamp 1018054153
transform 1 0 912 0 1 340
box -16 -6 32 210
use FILL  FILL_1309
timestamp 1018054153
transform 1 0 896 0 1 340
box -16 -6 32 210
use FILL  FILL_1310
timestamp 1018054153
transform 1 0 880 0 1 340
box -16 -6 32 210
use FILL  FILL_1311
timestamp 1018054153
transform 1 0 864 0 1 340
box -16 -6 32 210
use FILL  FILL_1312
timestamp 1018054153
transform 1 0 848 0 1 340
box -16 -6 32 210
use FILL  FILL_1313
timestamp 1018054153
transform 1 0 640 0 1 340
box -16 -6 32 210
use FILL  FILL_1314
timestamp 1018054153
transform 1 0 624 0 1 340
box -16 -6 32 210
use FILL  FILL_1315
timestamp 1018054153
transform 1 0 608 0 1 340
box -16 -6 32 210
use FILL  FILL_1316
timestamp 1018054153
transform 1 0 592 0 1 340
box -16 -6 32 210
use FILL  FILL_1317
timestamp 1018054153
transform 1 0 576 0 1 340
box -16 -6 32 210
use FILL  FILL_1318
timestamp 1018054153
transform 1 0 560 0 1 340
box -16 -6 32 210
use FILL  FILL_1319
timestamp 1018054153
transform 1 0 544 0 1 340
box -16 -6 32 210
use FILL  FILL_1320
timestamp 1018054153
transform 1 0 528 0 1 340
box -16 -6 32 210
use FILL  FILL_1321
timestamp 1018054153
transform 1 0 512 0 1 340
box -16 -6 32 210
use FILL  FILL_1322
timestamp 1018054153
transform 1 0 496 0 1 340
box -16 -6 32 210
use FILL  FILL_1323
timestamp 1018054153
transform 1 0 480 0 1 340
box -16 -6 32 210
use FILL  FILL_1324
timestamp 1018054153
transform 1 0 464 0 1 340
box -16 -6 32 210
use FILL  FILL_1325
timestamp 1018054153
transform 1 0 448 0 1 340
box -16 -6 32 210
use FILL  FILL_1326
timestamp 1018054153
transform 1 0 432 0 1 340
box -16 -6 32 210
use FILL  FILL_1327
timestamp 1018054153
transform 1 0 416 0 1 340
box -16 -6 32 210
use FILL  FILL_1328
timestamp 1018054153
transform 1 0 400 0 1 340
box -16 -6 32 210
use FILL  FILL_1329
timestamp 1018054153
transform 1 0 384 0 1 340
box -16 -6 32 210
use FILL  FILL_1330
timestamp 1018054153
transform 1 0 368 0 1 340
box -16 -6 32 210
use FILL  FILL_1331
timestamp 1018054153
transform 1 0 352 0 1 340
box -16 -6 32 210
use FILL  FILL_1332
timestamp 1018054153
transform 1 0 336 0 1 340
box -16 -6 32 210
use FILL  FILL_1333
timestamp 1018054153
transform 1 0 320 0 1 340
box -16 -6 32 210
use FILL  FILL_1334
timestamp 1018054153
transform 1 0 304 0 1 340
box -16 -6 32 210
use FILL  FILL_1335
timestamp 1018054153
transform 1 0 288 0 1 340
box -16 -6 32 210
use FILL  FILL_1336
timestamp 1018054153
transform 1 0 272 0 1 340
box -16 -6 32 210
use FILL  FILL_1337
timestamp 1018054153
transform 1 0 256 0 1 340
box -16 -6 32 210
use FILL  FILL_1338
timestamp 1018054153
transform 1 0 240 0 1 340
box -16 -6 32 210
use FILL  FILL_1339
timestamp 1018054153
transform 1 0 224 0 1 340
box -16 -6 32 210
use FILL  FILL_1340
timestamp 1018054153
transform 1 0 208 0 1 340
box -16 -6 32 210
use FILL  FILL_1341
timestamp 1018054153
transform 1 0 192 0 1 340
box -16 -6 32 210
use FILL  FILL_1342
timestamp 1018054153
transform 1 0 176 0 1 340
box -16 -6 32 210
use FILL  FILL_1343
timestamp 1018054153
transform 1 0 160 0 1 340
box -16 -6 32 210
use FILL  FILL_1344
timestamp 1018054153
transform 1 0 144 0 1 340
box -16 -6 32 210
use FILL  FILL_1345
timestamp 1018054153
transform 1 0 3664 0 -1 340
box -16 -6 32 210
use FILL  FILL_1346
timestamp 1018054153
transform 1 0 3648 0 -1 340
box -16 -6 32 210
use FILL  FILL_1347
timestamp 1018054153
transform 1 0 3632 0 -1 340
box -16 -6 32 210
use FILL  FILL_1348
timestamp 1018054153
transform 1 0 3616 0 -1 340
box -16 -6 32 210
use FILL  FILL_1349
timestamp 1018054153
transform 1 0 3600 0 -1 340
box -16 -6 32 210
use FILL  FILL_1350
timestamp 1018054153
transform 1 0 3584 0 -1 340
box -16 -6 32 210
use FILL  FILL_1351
timestamp 1018054153
transform 1 0 3568 0 -1 340
box -16 -6 32 210
use FILL  FILL_1352
timestamp 1018054153
transform 1 0 3552 0 -1 340
box -16 -6 32 210
use FILL  FILL_1353
timestamp 1018054153
transform 1 0 3536 0 -1 340
box -16 -6 32 210
use FILL  FILL_1354
timestamp 1018054153
transform 1 0 3520 0 -1 340
box -16 -6 32 210
use FILL  FILL_1355
timestamp 1018054153
transform 1 0 3504 0 -1 340
box -16 -6 32 210
use FILL  FILL_1356
timestamp 1018054153
transform 1 0 3488 0 -1 340
box -16 -6 32 210
use FILL  FILL_1357
timestamp 1018054153
transform 1 0 3472 0 -1 340
box -16 -6 32 210
use FILL  FILL_1358
timestamp 1018054153
transform 1 0 3456 0 -1 340
box -16 -6 32 210
use FILL  FILL_1359
timestamp 1018054153
transform 1 0 3440 0 -1 340
box -16 -6 32 210
use FILL  FILL_1360
timestamp 1018054153
transform 1 0 3424 0 -1 340
box -16 -6 32 210
use FILL  FILL_1361
timestamp 1018054153
transform 1 0 3408 0 -1 340
box -16 -6 32 210
use FILL  FILL_1362
timestamp 1018054153
transform 1 0 3392 0 -1 340
box -16 -6 32 210
use FILL  FILL_1363
timestamp 1018054153
transform 1 0 3376 0 -1 340
box -16 -6 32 210
use FILL  FILL_1364
timestamp 1018054153
transform 1 0 3360 0 -1 340
box -16 -6 32 210
use FILL  FILL_1365
timestamp 1018054153
transform 1 0 3344 0 -1 340
box -16 -6 32 210
use FILL  FILL_1366
timestamp 1018054153
transform 1 0 3328 0 -1 340
box -16 -6 32 210
use FILL  FILL_1367
timestamp 1018054153
transform 1 0 3312 0 -1 340
box -16 -6 32 210
use FILL  FILL_1368
timestamp 1018054153
transform 1 0 3296 0 -1 340
box -16 -6 32 210
use FILL  FILL_1369
timestamp 1018054153
transform 1 0 3280 0 -1 340
box -16 -6 32 210
use FILL  FILL_1370
timestamp 1018054153
transform 1 0 3264 0 -1 340
box -16 -6 32 210
use FILL  FILL_1371
timestamp 1018054153
transform 1 0 3248 0 -1 340
box -16 -6 32 210
use FILL  FILL_1372
timestamp 1018054153
transform 1 0 3200 0 -1 340
box -16 -6 32 210
use FILL  FILL_1373
timestamp 1018054153
transform 1 0 3184 0 -1 340
box -16 -6 32 210
use FILL  FILL_1374
timestamp 1018054153
transform 1 0 3168 0 -1 340
box -16 -6 32 210
use FILL  FILL_1375
timestamp 1018054153
transform 1 0 3152 0 -1 340
box -16 -6 32 210
use FILL  FILL_1376
timestamp 1018054153
transform 1 0 3136 0 -1 340
box -16 -6 32 210
use FILL  FILL_1377
timestamp 1018054153
transform 1 0 3120 0 -1 340
box -16 -6 32 210
use FILL  FILL_1378
timestamp 1018054153
transform 1 0 3104 0 -1 340
box -16 -6 32 210
use FILL  FILL_1379
timestamp 1018054153
transform 1 0 3088 0 -1 340
box -16 -6 32 210
use FILL  FILL_1380
timestamp 1018054153
transform 1 0 3072 0 -1 340
box -16 -6 32 210
use FILL  FILL_1381
timestamp 1018054153
transform 1 0 3008 0 -1 340
box -16 -6 32 210
use FILL  FILL_1382
timestamp 1018054153
transform 1 0 2992 0 -1 340
box -16 -6 32 210
use FILL  FILL_1383
timestamp 1018054153
transform 1 0 2976 0 -1 340
box -16 -6 32 210
use FILL  FILL_1384
timestamp 1018054153
transform 1 0 2832 0 -1 340
box -16 -6 32 210
use FILL  FILL_1385
timestamp 1018054153
transform 1 0 2608 0 -1 340
box -16 -6 32 210
use FILL  FILL_1386
timestamp 1018054153
transform 1 0 2592 0 -1 340
box -16 -6 32 210
use FILL  FILL_1387
timestamp 1018054153
transform 1 0 2576 0 -1 340
box -16 -6 32 210
use FILL  FILL_1388
timestamp 1018054153
transform 1 0 2560 0 -1 340
box -16 -6 32 210
use FILL  FILL_1389
timestamp 1018054153
transform 1 0 2512 0 -1 340
box -16 -6 32 210
use FILL  FILL_1390
timestamp 1018054153
transform 1 0 2496 0 -1 340
box -16 -6 32 210
use FILL  FILL_1391
timestamp 1018054153
transform 1 0 2480 0 -1 340
box -16 -6 32 210
use FILL  FILL_1392
timestamp 1018054153
transform 1 0 2464 0 -1 340
box -16 -6 32 210
use FILL  FILL_1393
timestamp 1018054153
transform 1 0 2448 0 -1 340
box -16 -6 32 210
use FILL  FILL_1394
timestamp 1018054153
transform 1 0 2432 0 -1 340
box -16 -6 32 210
use FILL  FILL_1395
timestamp 1018054153
transform 1 0 2416 0 -1 340
box -16 -6 32 210
use FILL  FILL_1396
timestamp 1018054153
transform 1 0 2400 0 -1 340
box -16 -6 32 210
use FILL  FILL_1397
timestamp 1018054153
transform 1 0 2384 0 -1 340
box -16 -6 32 210
use FILL  FILL_1398
timestamp 1018054153
transform 1 0 2368 0 -1 340
box -16 -6 32 210
use FILL  FILL_1399
timestamp 1018054153
transform 1 0 2352 0 -1 340
box -16 -6 32 210
use FILL  FILL_1400
timestamp 1018054153
transform 1 0 2336 0 -1 340
box -16 -6 32 210
use FILL  FILL_1401
timestamp 1018054153
transform 1 0 2320 0 -1 340
box -16 -6 32 210
use FILL  FILL_1402
timestamp 1018054153
transform 1 0 2304 0 -1 340
box -16 -6 32 210
use FILL  FILL_1403
timestamp 1018054153
transform 1 0 2288 0 -1 340
box -16 -6 32 210
use FILL  FILL_1404
timestamp 1018054153
transform 1 0 2272 0 -1 340
box -16 -6 32 210
use FILL  FILL_1405
timestamp 1018054153
transform 1 0 2256 0 -1 340
box -16 -6 32 210
use FILL  FILL_1406
timestamp 1018054153
transform 1 0 2240 0 -1 340
box -16 -6 32 210
use FILL  FILL_1407
timestamp 1018054153
transform 1 0 2224 0 -1 340
box -16 -6 32 210
use FILL  FILL_1408
timestamp 1018054153
transform 1 0 2208 0 -1 340
box -16 -6 32 210
use FILL  FILL_1409
timestamp 1018054153
transform 1 0 2192 0 -1 340
box -16 -6 32 210
use FILL  FILL_1410
timestamp 1018054153
transform 1 0 2176 0 -1 340
box -16 -6 32 210
use FILL  FILL_1411
timestamp 1018054153
transform 1 0 2160 0 -1 340
box -16 -6 32 210
use FILL  FILL_1412
timestamp 1018054153
transform 1 0 2144 0 -1 340
box -16 -6 32 210
use FILL  FILL_1413
timestamp 1018054153
transform 1 0 2128 0 -1 340
box -16 -6 32 210
use FILL  FILL_1414
timestamp 1018054153
transform 1 0 2112 0 -1 340
box -16 -6 32 210
use FILL  FILL_1415
timestamp 1018054153
transform 1 0 2096 0 -1 340
box -16 -6 32 210
use FILL  FILL_1416
timestamp 1018054153
transform 1 0 2080 0 -1 340
box -16 -6 32 210
use FILL  FILL_1417
timestamp 1018054153
transform 1 0 2064 0 -1 340
box -16 -6 32 210
use FILL  FILL_1418
timestamp 1018054153
transform 1 0 2048 0 -1 340
box -16 -6 32 210
use FILL  FILL_1419
timestamp 1018054153
transform 1 0 2032 0 -1 340
box -16 -6 32 210
use FILL  FILL_1420
timestamp 1018054153
transform 1 0 2016 0 -1 340
box -16 -6 32 210
use FILL  FILL_1421
timestamp 1018054153
transform 1 0 2000 0 -1 340
box -16 -6 32 210
use FILL  FILL_1422
timestamp 1018054153
transform 1 0 1984 0 -1 340
box -16 -6 32 210
use FILL  FILL_1423
timestamp 1018054153
transform 1 0 1968 0 -1 340
box -16 -6 32 210
use FILL  FILL_1424
timestamp 1018054153
transform 1 0 1952 0 -1 340
box -16 -6 32 210
use FILL  FILL_1425
timestamp 1018054153
transform 1 0 1936 0 -1 340
box -16 -6 32 210
use FILL  FILL_1426
timestamp 1018054153
transform 1 0 1920 0 -1 340
box -16 -6 32 210
use FILL  FILL_1427
timestamp 1018054153
transform 1 0 1904 0 -1 340
box -16 -6 32 210
use FILL  FILL_1428
timestamp 1018054153
transform 1 0 1888 0 -1 340
box -16 -6 32 210
use FILL  FILL_1429
timestamp 1018054153
transform 1 0 1872 0 -1 340
box -16 -6 32 210
use FILL  FILL_1430
timestamp 1018054153
transform 1 0 1856 0 -1 340
box -16 -6 32 210
use FILL  FILL_1431
timestamp 1018054153
transform 1 0 1840 0 -1 340
box -16 -6 32 210
use FILL  FILL_1432
timestamp 1018054153
transform 1 0 1824 0 -1 340
box -16 -6 32 210
use FILL  FILL_1433
timestamp 1018054153
transform 1 0 1808 0 -1 340
box -16 -6 32 210
use FILL  FILL_1434
timestamp 1018054153
transform 1 0 1792 0 -1 340
box -16 -6 32 210
use FILL  FILL_1435
timestamp 1018054153
transform 1 0 1776 0 -1 340
box -16 -6 32 210
use FILL  FILL_1436
timestamp 1018054153
transform 1 0 1664 0 -1 340
box -16 -6 32 210
use FILL  FILL_1437
timestamp 1018054153
transform 1 0 1648 0 -1 340
box -16 -6 32 210
use FILL  FILL_1438
timestamp 1018054153
transform 1 0 1632 0 -1 340
box -16 -6 32 210
use FILL  FILL_1439
timestamp 1018054153
transform 1 0 1616 0 -1 340
box -16 -6 32 210
use FILL  FILL_1440
timestamp 1018054153
transform 1 0 1600 0 -1 340
box -16 -6 32 210
use FILL  FILL_1441
timestamp 1018054153
transform 1 0 1536 0 -1 340
box -16 -6 32 210
use FILL  FILL_1442
timestamp 1018054153
transform 1 0 1520 0 -1 340
box -16 -6 32 210
use FILL  FILL_1443
timestamp 1018054153
transform 1 0 1440 0 -1 340
box -16 -6 32 210
use FILL  FILL_1444
timestamp 1018054153
transform 1 0 1424 0 -1 340
box -16 -6 32 210
use FILL  FILL_1445
timestamp 1018054153
transform 1 0 1408 0 -1 340
box -16 -6 32 210
use FILL  FILL_1446
timestamp 1018054153
transform 1 0 1392 0 -1 340
box -16 -6 32 210
use FILL  FILL_1447
timestamp 1018054153
transform 1 0 1376 0 -1 340
box -16 -6 32 210
use FILL  FILL_1448
timestamp 1018054153
transform 1 0 1360 0 -1 340
box -16 -6 32 210
use FILL  FILL_1449
timestamp 1018054153
transform 1 0 1120 0 -1 340
box -16 -6 32 210
use FILL  FILL_1450
timestamp 1018054153
transform 1 0 1104 0 -1 340
box -16 -6 32 210
use FILL  FILL_1451
timestamp 1018054153
transform 1 0 1088 0 -1 340
box -16 -6 32 210
use FILL  FILL_1452
timestamp 1018054153
transform 1 0 1072 0 -1 340
box -16 -6 32 210
use FILL  FILL_1453
timestamp 1018054153
transform 1 0 1056 0 -1 340
box -16 -6 32 210
use FILL  FILL_1454
timestamp 1018054153
transform 1 0 1040 0 -1 340
box -16 -6 32 210
use FILL  FILL_1455
timestamp 1018054153
transform 1 0 1024 0 -1 340
box -16 -6 32 210
use FILL  FILL_1456
timestamp 1018054153
transform 1 0 1008 0 -1 340
box -16 -6 32 210
use FILL  FILL_1457
timestamp 1018054153
transform 1 0 992 0 -1 340
box -16 -6 32 210
use FILL  FILL_1458
timestamp 1018054153
transform 1 0 976 0 -1 340
box -16 -6 32 210
use FILL  FILL_1459
timestamp 1018054153
transform 1 0 960 0 -1 340
box -16 -6 32 210
use FILL  FILL_1460
timestamp 1018054153
transform 1 0 944 0 -1 340
box -16 -6 32 210
use FILL  FILL_1461
timestamp 1018054153
transform 1 0 928 0 -1 340
box -16 -6 32 210
use FILL  FILL_1462
timestamp 1018054153
transform 1 0 912 0 -1 340
box -16 -6 32 210
use FILL  FILL_1463
timestamp 1018054153
transform 1 0 896 0 -1 340
box -16 -6 32 210
use FILL  FILL_1464
timestamp 1018054153
transform 1 0 880 0 -1 340
box -16 -6 32 210
use FILL  FILL_1465
timestamp 1018054153
transform 1 0 864 0 -1 340
box -16 -6 32 210
use FILL  FILL_1466
timestamp 1018054153
transform 1 0 848 0 -1 340
box -16 -6 32 210
use FILL  FILL_1467
timestamp 1018054153
transform 1 0 832 0 -1 340
box -16 -6 32 210
use FILL  FILL_1468
timestamp 1018054153
transform 1 0 816 0 -1 340
box -16 -6 32 210
use FILL  FILL_1469
timestamp 1018054153
transform 1 0 800 0 -1 340
box -16 -6 32 210
use FILL  FILL_1470
timestamp 1018054153
transform 1 0 784 0 -1 340
box -16 -6 32 210
use FILL  FILL_1471
timestamp 1018054153
transform 1 0 768 0 -1 340
box -16 -6 32 210
use FILL  FILL_1472
timestamp 1018054153
transform 1 0 752 0 -1 340
box -16 -6 32 210
use FILL  FILL_1473
timestamp 1018054153
transform 1 0 736 0 -1 340
box -16 -6 32 210
use FILL  FILL_1474
timestamp 1018054153
transform 1 0 720 0 -1 340
box -16 -6 32 210
use FILL  FILL_1475
timestamp 1018054153
transform 1 0 704 0 -1 340
box -16 -6 32 210
use FILL  FILL_1476
timestamp 1018054153
transform 1 0 688 0 -1 340
box -16 -6 32 210
use FILL  FILL_1477
timestamp 1018054153
transform 1 0 672 0 -1 340
box -16 -6 32 210
use FILL  FILL_1478
timestamp 1018054153
transform 1 0 656 0 -1 340
box -16 -6 32 210
use FILL  FILL_1479
timestamp 1018054153
transform 1 0 640 0 -1 340
box -16 -6 32 210
use FILL  FILL_1480
timestamp 1018054153
transform 1 0 624 0 -1 340
box -16 -6 32 210
use FILL  FILL_1481
timestamp 1018054153
transform 1 0 608 0 -1 340
box -16 -6 32 210
use FILL  FILL_1482
timestamp 1018054153
transform 1 0 592 0 -1 340
box -16 -6 32 210
use FILL  FILL_1483
timestamp 1018054153
transform 1 0 576 0 -1 340
box -16 -6 32 210
use FILL  FILL_1484
timestamp 1018054153
transform 1 0 560 0 -1 340
box -16 -6 32 210
use FILL  FILL_1485
timestamp 1018054153
transform 1 0 544 0 -1 340
box -16 -6 32 210
use FILL  FILL_1486
timestamp 1018054153
transform 1 0 528 0 -1 340
box -16 -6 32 210
use FILL  FILL_1487
timestamp 1018054153
transform 1 0 512 0 -1 340
box -16 -6 32 210
use FILL  FILL_1488
timestamp 1018054153
transform 1 0 496 0 -1 340
box -16 -6 32 210
use FILL  FILL_1489
timestamp 1018054153
transform 1 0 480 0 -1 340
box -16 -6 32 210
use FILL  FILL_1490
timestamp 1018054153
transform 1 0 464 0 -1 340
box -16 -6 32 210
use FILL  FILL_1491
timestamp 1018054153
transform 1 0 448 0 -1 340
box -16 -6 32 210
use FILL  FILL_1492
timestamp 1018054153
transform 1 0 432 0 -1 340
box -16 -6 32 210
use FILL  FILL_1493
timestamp 1018054153
transform 1 0 416 0 -1 340
box -16 -6 32 210
use FILL  FILL_1494
timestamp 1018054153
transform 1 0 400 0 -1 340
box -16 -6 32 210
use FILL  FILL_1495
timestamp 1018054153
transform 1 0 384 0 -1 340
box -16 -6 32 210
use FILL  FILL_1496
timestamp 1018054153
transform 1 0 368 0 -1 340
box -16 -6 32 210
use FILL  FILL_1497
timestamp 1018054153
transform 1 0 352 0 -1 340
box -16 -6 32 210
use FILL  FILL_1498
timestamp 1018054153
transform 1 0 336 0 -1 340
box -16 -6 32 210
use FILL  FILL_1499
timestamp 1018054153
transform 1 0 320 0 -1 340
box -16 -6 32 210
use FILL  FILL_1500
timestamp 1018054153
transform 1 0 304 0 -1 340
box -16 -6 32 210
use FILL  FILL_1501
timestamp 1018054153
transform 1 0 288 0 -1 340
box -16 -6 32 210
use FILL  FILL_1502
timestamp 1018054153
transform 1 0 272 0 -1 340
box -16 -6 32 210
use FILL  FILL_1503
timestamp 1018054153
transform 1 0 256 0 -1 340
box -16 -6 32 210
use FILL  FILL_1504
timestamp 1018054153
transform 1 0 240 0 -1 340
box -16 -6 32 210
use FILL  FILL_1505
timestamp 1018054153
transform 1 0 224 0 -1 340
box -16 -6 32 210
use FILL  FILL_1506
timestamp 1018054153
transform 1 0 208 0 -1 340
box -16 -6 32 210
use FILL  FILL_1507
timestamp 1018054153
transform 1 0 192 0 -1 340
box -16 -6 32 210
use FILL  FILL_1508
timestamp 1018054153
transform 1 0 176 0 -1 340
box -16 -6 32 210
use FILL  FILL_1509
timestamp 1018054153
transform 1 0 160 0 -1 340
box -16 -6 32 210
use FILL  FILL_1510
timestamp 1018054153
transform 1 0 144 0 -1 340
box -16 -6 32 210
use INVX1  INVX1_0
timestamp 1053022145
transform 1 0 3248 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_0
timestamp 1053022145
transform 1 0 3360 0 -1 1540
box -18 -6 52 210
use INVX2  INVX2_1
timestamp 1053022145
transform 1 0 3216 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_2
timestamp 1053022145
transform 1 0 3440 0 1 1140
box -18 -6 52 210
use INVX2  INVX2_3
timestamp 1053022145
transform 1 0 3488 0 -1 1540
box -18 -6 52 210
use INVX2  INVX2_4
timestamp 1053022145
transform 1 0 3360 0 -1 1140
box -18 -6 52 210
use INVX2  INVX2_5
timestamp 1053022145
transform 1 0 3568 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_6
timestamp 1053022145
transform 1 0 3360 0 1 740
box -18 -6 52 210
use INVX2  INVX2_7
timestamp 1053022145
transform 1 0 3344 0 1 340
box -18 -6 52 210
use INVX2  INVX2_8
timestamp 1053022145
transform 1 0 3072 0 1 340
box -18 -6 52 210
use INVX2  INVX2_9
timestamp 1053022145
transform 1 0 3216 0 -1 340
box -18 -6 52 210
use INVX2  INVX2_10
timestamp 1053022145
transform 1 0 2944 0 -1 340
box -18 -6 52 210
use INVX2  INVX2_11
timestamp 1053022145
transform 1 0 2624 0 1 340
box -18 -6 52 210
use INVX2  INVX2_12
timestamp 1053022145
transform 1 0 2528 0 -1 340
box -18 -6 52 210
use INVX2  INVX2_13
timestamp 1053022145
transform 1 0 2416 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_14
timestamp 1053022145
transform 1 0 2512 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_15
timestamp 1053022145
transform 1 0 2176 0 1 340
box -18 -6 52 210
use INVX2  INVX2_16
timestamp 1053022145
transform 1 0 2224 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_17
timestamp 1053022145
transform 1 0 2656 0 -1 1140
box -18 -6 52 210
use INVX2  INVX2_18
timestamp 1053022145
transform 1 0 2304 0 1 1140
box -18 -6 52 210
use INVX2  INVX2_19
timestamp 1053022145
transform 1 0 1296 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_20
timestamp 1053022145
transform 1 0 560 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_21
timestamp 1053022145
transform 1 0 944 0 -1 1540
box -18 -6 52 210
use INVX2  INVX2_22
timestamp 1053022145
transform 1 0 736 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_23
timestamp 1053022145
transform 1 0 512 0 1 1140
box -18 -6 52 210
use INVX2  INVX2_24
timestamp 1053022145
transform 1 0 2752 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_25
timestamp 1053022145
transform 1 0 2496 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_26
timestamp 1053022145
transform 1 0 1680 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_27
timestamp 1053022145
transform 1 0 1680 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_28
timestamp 1053022145
transform 1 0 1664 0 1 1140
box -18 -6 52 210
use INVX2  INVX2_29
timestamp 1053022145
transform 1 0 1776 0 -1 1140
box -18 -6 52 210
use INVX2  INVX2_30
timestamp 1053022145
transform 1 0 2176 0 -1 1140
box -18 -6 52 210
use INVX2  INVX2_31
timestamp 1053022145
transform 1 0 2288 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_32
timestamp 1053022145
transform 1 0 1552 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_33
timestamp 1053022145
transform 1 0 1152 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_34
timestamp 1053022145
transform 1 0 800 0 -1 1540
box -18 -6 52 210
use INVX2  INVX2_35
timestamp 1053022145
transform 1 0 2096 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_36
timestamp 1053022145
transform 1 0 2128 0 -1 2340
box -18 -6 52 210
use INVX2  INVX2_37
timestamp 1053022145
transform 1 0 1328 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_38
timestamp 1053022145
transform 1 0 1632 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_39
timestamp 1053022145
transform 1 0 2336 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_40
timestamp 1053022145
transform 1 0 3104 0 -1 2740
box -18 -6 52 210
use INVX2  INVX2_41
timestamp 1053022145
transform 1 0 864 0 -1 2740
box -18 -6 52 210
use INVX2  INVX2_42
timestamp 1053022145
transform 1 0 1008 0 1 2340
box -18 -6 52 210
use INVX2  INVX2_43
timestamp 1053022145
transform 1 0 3328 0 -1 2740
box -18 -6 52 210
use INVX2  INVX2_44
timestamp 1053022145
transform 1 0 512 0 1 2740
box -18 -6 52 210
use INVX2  INVX2_45
timestamp 1053022145
transform 1 0 2224 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_46
timestamp 1053022145
transform 1 0 2704 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_47
timestamp 1053022145
transform 1 0 3040 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_48
timestamp 1053022145
transform 1 0 2608 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_49
timestamp 1053022145
transform 1 0 656 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_50
timestamp 1053022145
transform 1 0 2928 0 -1 3140
box -18 -6 52 210
use INVX2  INVX2_51
timestamp 1053022145
transform 1 0 1024 0 -1 3140
box -18 -6 52 210
use INVX2  INVX2_52
timestamp 1053022145
transform 1 0 1248 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_53
timestamp 1053022145
transform 1 0 2992 0 1 2740
box -18 -6 52 210
use INVX2  INVX2_54
timestamp 1053022145
transform 1 0 1008 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_55
timestamp 1053022145
transform 1 0 2848 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_56
timestamp 1053022145
transform 1 0 784 0 -1 2340
box -18 -6 52 210
use INVX2  INVX2_57
timestamp 1053022145
transform 1 0 1216 0 -1 2340
box -18 -6 52 210
use INVX2  INVX2_58
timestamp 1053022145
transform 1 0 3248 0 -1 2340
box -18 -6 52 210
use INVX2  INVX2_59
timestamp 1053022145
transform 1 0 1696 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_60
timestamp 1053022145
transform 1 0 1472 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_61
timestamp 1053022145
transform 1 0 976 0 1 3140
box -18 -6 52 210
use INVX2  INVX2_62
timestamp 1053022145
transform 1 0 352 0 -1 3140
box -18 -6 52 210
use INVX2  INVX2_63
timestamp 1053022145
transform 1 0 1616 0 1 340
box -18 -6 52 210
use INVX2  INVX2_64
timestamp 1053022145
transform 1 0 1504 0 1 340
box -18 -6 52 210
use INVX2  INVX2_65
timestamp 1053022145
transform 1 0 560 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_66
timestamp 1053022145
transform 1 0 896 0 1 740
box -18 -6 52 210
use INVX2  INVX2_67
timestamp 1053022145
transform 1 0 2432 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_68
timestamp 1053022145
transform 1 0 1920 0 -1 1140
box -18 -6 52 210
use INVX2  INVX2_69
timestamp 1053022145
transform 1 0 1296 0 1 740
box -18 -6 52 210
use INVX2  INVX2_70
timestamp 1053022145
transform 1 0 1984 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_71
timestamp 1053022145
transform 1 0 1920 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_72
timestamp 1053022145
transform 1 0 816 0 1 1540
box -18 -6 52 210
use INVX2  INVX2_73
timestamp 1053022145
transform 1 0 1248 0 1 740
box -18 -6 52 210
use INVX2  INVX2_74
timestamp 1053022145
transform 1 0 768 0 1 740
box -18 -6 52 210
use INVX2  INVX2_75
timestamp 1053022145
transform 1 0 2720 0 1 1140
box -18 -6 52 210
use INVX2  INVX2_76
timestamp 1053022145
transform 1 0 2032 0 1 340
box -18 -6 52 210
use INVX2  INVX2_77
timestamp 1053022145
transform 1 0 2048 0 -1 740
box -18 -6 52 210
use INVX2  INVX2_78
timestamp 1053022145
transform 1 0 2352 0 1 740
box -18 -6 52 210
use INVX2  INVX2_79
timestamp 1053022145
transform 1 0 3344 0 1 2740
box -18 -6 52 210
use INVX2  INVX2_80
timestamp 1053022145
transform 1 0 576 0 1 2340
box -18 -6 52 210
use INVX2  INVX2_81
timestamp 1053022145
transform 1 0 528 0 -1 2740
box -18 -6 52 210
use INVX2  INVX2_82
timestamp 1053022145
transform 1 0 3072 0 1 2340
box -18 -6 52 210
use INVX2  INVX2_83
timestamp 1053022145
transform 1 0 2912 0 -1 2340
box -18 -6 52 210
use INVX2  INVX2_84
timestamp 1053022145
transform 1 0 832 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_85
timestamp 1053022145
transform 1 0 640 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_86
timestamp 1053022145
transform 1 0 3040 0 1 1940
box -18 -6 52 210
use INVX2  INVX2_87
timestamp 1053022145
transform 1 0 3104 0 1 2740
box -18 -6 52 210
use INVX2  INVX2_88
timestamp 1053022145
transform 1 0 1216 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_89
timestamp 1053022145
transform 1 0 720 0 -1 3140
box -18 -6 52 210
use INVX2  INVX2_90
timestamp 1053022145
transform 1 0 3280 0 -1 3140
box -18 -6 52 210
use INVX2  INVX2_91
timestamp 1053022145
transform 1 0 2448 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_92
timestamp 1053022145
transform 1 0 3216 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_93
timestamp 1053022145
transform 1 0 2864 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_94
timestamp 1053022145
transform 1 0 2192 0 -1 3540
box -18 -6 52 210
use INVX2  INVX2_95
timestamp 1053022145
transform 1 0 1744 0 -1 340
box -18 -6 52 210
use INVX2  INVX2_96
timestamp 1053022145
transform 1 0 1328 0 -1 340
box -18 -6 52 210
use INVX2  INVX2_97
timestamp 1053022145
transform 1 0 960 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_98
timestamp 1053022145
transform 1 0 928 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_99
timestamp 1053022145
transform 1 0 2224 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_100
timestamp 1053022145
transform 1 0 2256 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_101
timestamp 1053022145
transform 1 0 2288 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_102
timestamp 1053022145
transform 1 0 2880 0 -1 1940
box -18 -6 52 210
use INVX2  INVX2_103
timestamp 1053022145
transform 1 0 2576 0 1 740
box -18 -6 52 210
use INVX4  INVX4_0
timestamp 1053722803
transform 1 0 3200 0 1 1940
box -18 -6 56 210
use M2_M1  M2_M1_0
timestamp 1543120812
transform 1 0 2744 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_1
timestamp 1543120812
transform 1 0 2616 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_2
timestamp 1543120812
transform 1 0 2552 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_3
timestamp 1543120812
transform 1 0 2280 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_4
timestamp 1543120812
transform 1 0 2280 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_5
timestamp 1543120812
transform 1 0 3160 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_6
timestamp 1543120812
transform 1 0 2840 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_7
timestamp 1543120812
transform 1 0 2824 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_8
timestamp 1543120812
transform 1 0 2776 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_9
timestamp 1543120812
transform 1 0 2776 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_10
timestamp 1543120812
transform 1 0 2632 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_11
timestamp 1543120812
transform 1 0 3576 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_12
timestamp 1543120812
transform 1 0 3384 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_13
timestamp 1543120812
transform 1 0 3256 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_14
timestamp 1543120812
transform 1 0 3256 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_15
timestamp 1543120812
transform 1 0 3160 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_16
timestamp 1543120812
transform 1 0 3144 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_17
timestamp 1543120812
transform 1 0 3480 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_18
timestamp 1543120812
transform 1 0 3416 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_19
timestamp 1543120812
transform 1 0 3400 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_20
timestamp 1543120812
transform 1 0 3272 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_21
timestamp 1543120812
transform 1 0 3272 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_22
timestamp 1543120812
transform 1 0 3400 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_23
timestamp 1543120812
transform 1 0 3400 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_24
timestamp 1543120812
transform 1 0 3256 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_25
timestamp 1543120812
transform 1 0 3240 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_26
timestamp 1543120812
transform 1 0 3240 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_27
timestamp 1543120812
transform 1 0 2936 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_28
timestamp 1543120812
transform 1 0 2904 0 1 790
box -4 -4 4 4
use M2_M1  M2_M1_29
timestamp 1543120812
transform 1 0 2680 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_30
timestamp 1543120812
transform 1 0 2632 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_31
timestamp 1543120812
transform 1 0 2888 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_32
timestamp 1543120812
transform 1 0 2872 0 1 690
box -4 -4 4 4
use M2_M1  M2_M1_33
timestamp 1543120812
transform 1 0 2840 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_34
timestamp 1543120812
transform 1 0 2792 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_35
timestamp 1543120812
transform 1 0 3208 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_36
timestamp 1543120812
transform 1 0 3160 0 1 790
box -4 -4 4 4
use M2_M1  M2_M1_37
timestamp 1543120812
transform 1 0 3160 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_38
timestamp 1543120812
transform 1 0 3128 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_39
timestamp 1543120812
transform 1 0 3336 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_40
timestamp 1543120812
transform 1 0 3288 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_41
timestamp 1543120812
transform 1 0 3160 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_42
timestamp 1543120812
transform 1 0 3144 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_43
timestamp 1543120812
transform 1 0 3000 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_44
timestamp 1543120812
transform 1 0 3304 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_45
timestamp 1543120812
transform 1 0 3256 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_46
timestamp 1543120812
transform 1 0 3128 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_47
timestamp 1543120812
transform 1 0 3128 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_48
timestamp 1543120812
transform 1 0 3368 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_49
timestamp 1543120812
transform 1 0 3288 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_50
timestamp 1543120812
transform 1 0 3288 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_51
timestamp 1543120812
transform 1 0 3224 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_52
timestamp 1543120812
transform 1 0 3048 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_53
timestamp 1543120812
transform 1 0 3032 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_54
timestamp 1543120812
transform 1 0 3432 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_55
timestamp 1543120812
transform 1 0 3400 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_56
timestamp 1543120812
transform 1 0 3160 0 1 1590
box -4 -4 4 4
use M2_M1  M2_M1_57
timestamp 1543120812
transform 1 0 3096 0 1 1590
box -4 -4 4 4
use M2_M1  M2_M1_58
timestamp 1543120812
transform 1 0 3016 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_59
timestamp 1543120812
transform 1 0 3432 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_60
timestamp 1543120812
transform 1 0 3304 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_61
timestamp 1543120812
transform 1 0 3176 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_62
timestamp 1543120812
transform 1 0 2936 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_63
timestamp 1543120812
transform 1 0 2712 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_64
timestamp 1543120812
transform 1 0 2648 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_65
timestamp 1543120812
transform 1 0 2584 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_66
timestamp 1543120812
transform 1 0 2136 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_67
timestamp 1543120812
transform 1 0 2104 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_68
timestamp 1543120812
transform 1 0 1992 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_69
timestamp 1543120812
transform 1 0 2024 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_70
timestamp 1543120812
transform 1 0 2024 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_71
timestamp 1543120812
transform 1 0 1960 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_72
timestamp 1543120812
transform 1 0 1576 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_73
timestamp 1543120812
transform 1 0 1544 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_74
timestamp 1543120812
transform 1 0 1480 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_75
timestamp 1543120812
transform 1 0 1432 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_76
timestamp 1543120812
transform 1 0 2152 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_77
timestamp 1543120812
transform 1 0 2056 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_78
timestamp 1543120812
transform 1 0 1816 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_79
timestamp 1543120812
transform 1 0 1512 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_80
timestamp 1543120812
transform 1 0 1464 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_81
timestamp 1543120812
transform 1 0 1320 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_82
timestamp 1543120812
transform 1 0 2504 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_83
timestamp 1543120812
transform 1 0 2440 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_84
timestamp 1543120812
transform 1 0 2344 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_85
timestamp 1543120812
transform 1 0 2072 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_86
timestamp 1543120812
transform 1 0 2040 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_87
timestamp 1543120812
transform 1 0 2024 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_88
timestamp 1543120812
transform 1 0 1352 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_89
timestamp 1543120812
transform 1 0 1336 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_90
timestamp 1543120812
transform 1 0 1304 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_91
timestamp 1543120812
transform 1 0 1000 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_92
timestamp 1543120812
transform 1 0 984 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_93
timestamp 1543120812
transform 1 0 936 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_94
timestamp 1543120812
transform 1 0 840 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_95
timestamp 1543120812
transform 1 0 744 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_96
timestamp 1543120812
transform 1 0 936 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_97
timestamp 1543120812
transform 1 0 920 0 1 1270
box -4 -4 4 4
use M2_M1  M2_M1_98
timestamp 1543120812
transform 1 0 552 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_99
timestamp 1543120812
transform 1 0 520 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_100
timestamp 1543120812
transform 1 0 504 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_101
timestamp 1543120812
transform 1 0 1112 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_102
timestamp 1543120812
transform 1 0 1000 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_103
timestamp 1543120812
transform 1 0 680 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_104
timestamp 1543120812
transform 1 0 680 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_105
timestamp 1543120812
transform 1 0 552 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_106
timestamp 1543120812
transform 1 0 520 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_107
timestamp 1543120812
transform 1 0 2920 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_108
timestamp 1543120812
transform 1 0 2904 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_109
timestamp 1543120812
transform 1 0 2904 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_110
timestamp 1543120812
transform 1 0 2760 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_111
timestamp 1543120812
transform 1 0 2744 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_112
timestamp 1543120812
transform 1 0 1736 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_113
timestamp 1543120812
transform 1 0 1704 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_114
timestamp 1543120812
transform 1 0 1688 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_115
timestamp 1543120812
transform 1 0 1656 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_116
timestamp 1543120812
transform 1 0 1640 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_117
timestamp 1543120812
transform 1 0 1560 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_118
timestamp 1543120812
transform 1 0 1976 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_119
timestamp 1543120812
transform 1 0 1912 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_120
timestamp 1543120812
transform 1 0 1848 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_121
timestamp 1543120812
transform 1 0 1736 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_122
timestamp 1543120812
transform 1 0 1688 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_123
timestamp 1543120812
transform 1 0 1464 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_124
timestamp 1543120812
transform 1 0 1448 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_125
timestamp 1543120812
transform 1 0 2808 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_126
timestamp 1543120812
transform 1 0 2808 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_127
timestamp 1543120812
transform 1 0 2776 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_128
timestamp 1543120812
transform 1 0 2744 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_129
timestamp 1543120812
transform 1 0 2504 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_130
timestamp 1543120812
transform 1 0 2360 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_131
timestamp 1543120812
transform 1 0 2632 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_132
timestamp 1543120812
transform 1 0 2616 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_133
timestamp 1543120812
transform 1 0 2520 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_134
timestamp 1543120812
transform 1 0 2376 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_135
timestamp 1543120812
transform 1 0 2360 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_136
timestamp 1543120812
transform 1 0 2312 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_137
timestamp 1543120812
transform 1 0 1960 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_138
timestamp 1543120812
transform 1 0 1832 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_139
timestamp 1543120812
transform 1 0 1768 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_140
timestamp 1543120812
transform 1 0 1576 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_141
timestamp 1543120812
transform 1 0 1528 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_142
timestamp 1543120812
transform 1 0 1432 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_143
timestamp 1543120812
transform 1 0 1336 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_144
timestamp 1543120812
transform 1 0 1880 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_145
timestamp 1543120812
transform 1 0 1848 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_146
timestamp 1543120812
transform 1 0 1784 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_147
timestamp 1543120812
transform 1 0 1720 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_148
timestamp 1543120812
transform 1 0 1672 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_149
timestamp 1543120812
transform 1 0 1608 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_150
timestamp 1543120812
transform 1 0 1224 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_151
timestamp 1543120812
transform 1 0 2520 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_152
timestamp 1543120812
transform 1 0 2472 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_153
timestamp 1543120812
transform 1 0 2472 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_154
timestamp 1543120812
transform 1 0 2216 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_155
timestamp 1543120812
transform 1 0 2200 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_156
timestamp 1543120812
transform 1 0 2184 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_157
timestamp 1543120812
transform 1 0 2648 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_158
timestamp 1543120812
transform 1 0 2632 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_159
timestamp 1543120812
transform 1 0 2472 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_160
timestamp 1543120812
transform 1 0 2424 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_161
timestamp 1543120812
transform 1 0 2408 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_162
timestamp 1543120812
transform 1 0 2296 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_163
timestamp 1543120812
transform 1 0 2232 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_164
timestamp 1543120812
transform 1 0 1576 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_165
timestamp 1543120812
transform 1 0 1560 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_166
timestamp 1543120812
transform 1 0 1496 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_167
timestamp 1543120812
transform 1 0 1464 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_168
timestamp 1543120812
transform 1 0 1304 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_169
timestamp 1543120812
transform 1 0 1208 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_170
timestamp 1543120812
transform 1 0 1176 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_171
timestamp 1543120812
transform 1 0 1464 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_172
timestamp 1543120812
transform 1 0 1416 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_173
timestamp 1543120812
transform 1 0 1336 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_174
timestamp 1543120812
transform 1 0 1224 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_175
timestamp 1543120812
transform 1 0 1160 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_176
timestamp 1543120812
transform 1 0 984 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_177
timestamp 1543120812
transform 1 0 952 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_178
timestamp 1543120812
transform 1 0 2520 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_179
timestamp 1543120812
transform 1 0 2488 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_180
timestamp 1543120812
transform 1 0 2136 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_181
timestamp 1543120812
transform 1 0 2120 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_182
timestamp 1543120812
transform 1 0 2104 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_183
timestamp 1543120812
transform 1 0 2088 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_184
timestamp 1543120812
transform 1 0 2024 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_185
timestamp 1543120812
transform 1 0 2696 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_186
timestamp 1543120812
transform 1 0 2632 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_187
timestamp 1543120812
transform 1 0 2360 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_188
timestamp 1543120812
transform 1 0 2328 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_189
timestamp 1543120812
transform 1 0 2200 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_190
timestamp 1543120812
transform 1 0 1640 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_191
timestamp 1543120812
transform 1 0 1544 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_192
timestamp 1543120812
transform 1 0 1528 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_193
timestamp 1543120812
transform 1 0 1512 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_194
timestamp 1543120812
transform 1 0 1176 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_195
timestamp 1543120812
transform 1 0 1048 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_196
timestamp 1543120812
transform 1 0 1400 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_197
timestamp 1543120812
transform 1 0 1336 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_198
timestamp 1543120812
transform 1 0 1320 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_199
timestamp 1543120812
transform 1 0 1256 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_200
timestamp 1543120812
transform 1 0 1064 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_201
timestamp 1543120812
transform 1 0 904 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_202
timestamp 1543120812
transform 1 0 2744 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_203
timestamp 1543120812
transform 1 0 2504 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_204
timestamp 1543120812
transform 1 0 2200 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_205
timestamp 1543120812
transform 1 0 2136 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_206
timestamp 1543120812
transform 1 0 2120 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_207
timestamp 1543120812
transform 1 0 2040 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_208
timestamp 1543120812
transform 1 0 2616 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_209
timestamp 1543120812
transform 1 0 2312 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_210
timestamp 1543120812
transform 1 0 2264 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_211
timestamp 1543120812
transform 1 0 3160 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_212
timestamp 1543120812
transform 1 0 2904 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_213
timestamp 1543120812
transform 1 0 1736 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_214
timestamp 1543120812
transform 1 0 1624 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_215
timestamp 1543120812
transform 1 0 1544 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_216
timestamp 1543120812
transform 1 0 1400 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_217
timestamp 1543120812
transform 1 0 2936 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_218
timestamp 1543120812
transform 1 0 2712 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_219
timestamp 1543120812
transform 1 0 1624 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_220
timestamp 1543120812
transform 1 0 1352 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_221
timestamp 1543120812
transform 1 0 1336 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_222
timestamp 1543120812
transform 1 0 2232 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_223
timestamp 1543120812
transform 1 0 2136 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_224
timestamp 1543120812
transform 1 0 2104 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_225
timestamp 1543120812
transform 1 0 1928 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_226
timestamp 1543120812
transform 1 0 3000 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_227
timestamp 1543120812
transform 1 0 2984 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_228
timestamp 1543120812
transform 1 0 2824 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_229
timestamp 1543120812
transform 1 0 1464 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_230
timestamp 1543120812
transform 1 0 1240 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_231
timestamp 1543120812
transform 1 0 1240 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_232
timestamp 1543120812
transform 1 0 1352 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_233
timestamp 1543120812
transform 1 0 1128 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_234
timestamp 1543120812
transform 1 0 1032 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_235
timestamp 1543120812
transform 1 0 3144 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_236
timestamp 1543120812
transform 1 0 2936 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_237
timestamp 1543120812
transform 1 0 2712 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_238
timestamp 1543120812
transform 1 0 1224 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_239
timestamp 1543120812
transform 1 0 1128 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_240
timestamp 1543120812
transform 1 0 1112 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_241
timestamp 1543120812
transform 1 0 824 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_242
timestamp 1543120812
transform 1 0 792 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_243
timestamp 1543120812
transform 1 0 1144 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_244
timestamp 1543120812
transform 1 0 984 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_245
timestamp 1543120812
transform 1 0 968 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_246
timestamp 1543120812
transform 1 0 1000 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_247
timestamp 1543120812
transform 1 0 872 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_248
timestamp 1543120812
transform 1 0 2760 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_249
timestamp 1543120812
transform 1 0 2664 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_250
timestamp 1543120812
transform 1 0 2616 0 1 390
box -4 -4 4 4
use M2_M1  M2_M1_251
timestamp 1543120812
transform 1 0 3112 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_252
timestamp 1543120812
transform 1 0 3048 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_253
timestamp 1543120812
transform 1 0 3048 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_254
timestamp 1543120812
transform 1 0 3672 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_255
timestamp 1543120812
transform 1 0 3400 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_256
timestamp 1543120812
transform 1 0 3368 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_257
timestamp 1543120812
transform 1 0 3400 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_258
timestamp 1543120812
transform 1 0 3256 0 1 1890
box -4 -4 4 4
use M2_M1  M2_M1_259
timestamp 1543120812
transform 1 0 3208 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_260
timestamp 1543120812
transform 1 0 3496 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_261
timestamp 1543120812
transform 1 0 3432 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_262
timestamp 1543120812
transform 1 0 3480 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_263
timestamp 1543120812
transform 1 0 3448 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_264
timestamp 1543120812
transform 1 0 3384 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_265
timestamp 1543120812
transform 1 0 3400 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_266
timestamp 1543120812
transform 1 0 3352 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_267
timestamp 1543120812
transform 1 0 3336 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_268
timestamp 1543120812
transform 1 0 3320 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_269
timestamp 1543120812
transform 1 0 3560 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_270
timestamp 1543120812
transform 1 0 3544 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_271
timestamp 1543120812
transform 1 0 3576 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_272
timestamp 1543120812
transform 1 0 3576 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_273
timestamp 1543120812
transform 1 0 3528 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_274
timestamp 1543120812
transform 1 0 3368 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_275
timestamp 1543120812
transform 1 0 3336 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_276
timestamp 1543120812
transform 1 0 3352 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_277
timestamp 1543120812
transform 1 0 3352 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_278
timestamp 1543120812
transform 1 0 3320 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_279
timestamp 1543120812
transform 1 0 3320 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_280
timestamp 1543120812
transform 1 0 3240 0 1 450
box -4 -4 4 4
use M2_M1  M2_M1_281
timestamp 1543120812
transform 1 0 3496 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_282
timestamp 1543120812
transform 1 0 3112 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_283
timestamp 1543120812
transform 1 0 3080 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_284
timestamp 1543120812
transform 1 0 3320 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_285
timestamp 1543120812
transform 1 0 3224 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_286
timestamp 1543120812
transform 1 0 3224 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_287
timestamp 1543120812
transform 1 0 2952 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_288
timestamp 1543120812
transform 1 0 2888 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_289
timestamp 1543120812
transform 1 0 2808 0 1 450
box -4 -4 4 4
use M2_M1  M2_M1_290
timestamp 1543120812
transform 1 0 2696 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_291
timestamp 1543120812
transform 1 0 2664 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_292
timestamp 1543120812
transform 1 0 2632 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_293
timestamp 1543120812
transform 1 0 2920 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_294
timestamp 1543120812
transform 1 0 2536 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_295
timestamp 1543120812
transform 1 0 2840 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_296
timestamp 1543120812
transform 1 0 2424 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_297
timestamp 1543120812
transform 1 0 2392 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_298
timestamp 1543120812
transform 1 0 2616 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_299
timestamp 1543120812
transform 1 0 2504 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_300
timestamp 1543120812
transform 1 0 2344 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_301
timestamp 1543120812
transform 1 0 2184 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_302
timestamp 1543120812
transform 1 0 2392 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_303
timestamp 1543120812
transform 1 0 2232 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_304
timestamp 1543120812
transform 1 0 2696 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_305
timestamp 1543120812
transform 1 0 2664 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_306
timestamp 1543120812
transform 1 0 3288 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_307
timestamp 1543120812
transform 1 0 3256 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_308
timestamp 1543120812
transform 1 0 3560 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_309
timestamp 1543120812
transform 1 0 3496 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_310
timestamp 1543120812
transform 1 0 3448 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_311
timestamp 1543120812
transform 1 0 3608 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_312
timestamp 1543120812
transform 1 0 3512 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_313
timestamp 1543120812
transform 1 0 3512 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_314
timestamp 1543120812
transform 1 0 3464 0 1 1090
box -4 -4 4 4
use M2_M1  M2_M1_315
timestamp 1543120812
transform 1 0 3496 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_316
timestamp 1543120812
transform 1 0 3464 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_317
timestamp 1543120812
transform 1 0 3384 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_318
timestamp 1543120812
transform 1 0 3288 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_319
timestamp 1543120812
transform 1 0 3592 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_320
timestamp 1543120812
transform 1 0 3336 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_321
timestamp 1543120812
transform 1 0 3272 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_322
timestamp 1543120812
transform 1 0 3624 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_323
timestamp 1543120812
transform 1 0 3464 0 1 690
box -4 -4 4 4
use M2_M1  M2_M1_324
timestamp 1543120812
transform 1 0 3448 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_325
timestamp 1543120812
transform 1 0 3384 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_326
timestamp 1543120812
transform 1 0 3512 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_327
timestamp 1543120812
transform 1 0 3512 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_328
timestamp 1543120812
transform 1 0 3336 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_329
timestamp 1543120812
transform 1 0 3272 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_330
timestamp 1543120812
transform 1 0 3016 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_331
timestamp 1543120812
transform 1 0 2904 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_332
timestamp 1543120812
transform 1 0 2840 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_333
timestamp 1543120812
transform 1 0 3080 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_334
timestamp 1543120812
transform 1 0 2984 0 1 290
box -4 -4 4 4
use M2_M1  M2_M1_335
timestamp 1543120812
transform 1 0 2824 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_336
timestamp 1543120812
transform 1 0 2648 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_337
timestamp 1543120812
transform 1 0 3064 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_338
timestamp 1543120812
transform 1 0 2968 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_339
timestamp 1543120812
transform 1 0 2872 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_340
timestamp 1543120812
transform 1 0 2728 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_341
timestamp 1543120812
transform 1 0 2632 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_342
timestamp 1543120812
transform 1 0 2568 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_343
timestamp 1543120812
transform 1 0 2568 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_344
timestamp 1543120812
transform 1 0 2504 0 1 390
box -4 -4 4 4
use M2_M1  M2_M1_345
timestamp 1543120812
transform 1 0 2504 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_346
timestamp 1543120812
transform 1 0 2296 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_347
timestamp 1543120812
transform 1 0 2296 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_348
timestamp 1543120812
transform 1 0 2536 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_349
timestamp 1543120812
transform 1 0 2408 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_350
timestamp 1543120812
transform 1 0 2360 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_351
timestamp 1543120812
transform 1 0 2344 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_352
timestamp 1543120812
transform 1 0 2488 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_353
timestamp 1543120812
transform 1 0 2440 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_354
timestamp 1543120812
transform 1 0 2088 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_355
timestamp 1543120812
transform 1 0 2088 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_356
timestamp 1543120812
transform 1 0 2168 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_357
timestamp 1543120812
transform 1 0 1896 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_358
timestamp 1543120812
transform 1 0 2664 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_359
timestamp 1543120812
transform 1 0 2584 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_360
timestamp 1543120812
transform 1 0 2296 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_361
timestamp 1543120812
transform 1 0 2136 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_362
timestamp 1543120812
transform 1 0 2088 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_363
timestamp 1543120812
transform 1 0 1224 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_364
timestamp 1543120812
transform 1 0 1224 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_365
timestamp 1543120812
transform 1 0 1192 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_366
timestamp 1543120812
transform 1 0 1128 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_367
timestamp 1543120812
transform 1 0 1128 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_368
timestamp 1543120812
transform 1 0 952 0 1 690
box -4 -4 4 4
use M2_M1  M2_M1_369
timestamp 1543120812
transform 1 0 664 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_370
timestamp 1543120812
transform 1 0 632 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_371
timestamp 1543120812
transform 1 0 1048 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_372
timestamp 1543120812
transform 1 0 1016 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_373
timestamp 1543120812
transform 1 0 760 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_374
timestamp 1543120812
transform 1 0 632 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_375
timestamp 1543120812
transform 1 0 632 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_376
timestamp 1543120812
transform 1 0 552 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_377
timestamp 1543120812
transform 1 0 520 0 1 790
box -4 -4 4 4
use M2_M1  M2_M1_378
timestamp 1543120812
transform 1 0 1048 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_379
timestamp 1543120812
transform 1 0 1048 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_380
timestamp 1543120812
transform 1 0 520 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_381
timestamp 1543120812
transform 1 0 488 0 1 1490
box -4 -4 4 4
use M2_M1  M2_M1_382
timestamp 1543120812
transform 1 0 488 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_383
timestamp 1543120812
transform 1 0 2776 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_384
timestamp 1543120812
transform 1 0 2696 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_385
timestamp 1543120812
transform 1 0 2472 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_386
timestamp 1543120812
transform 1 0 2536 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_387
timestamp 1543120812
transform 1 0 2520 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_388
timestamp 1543120812
transform 1 0 2424 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_389
timestamp 1543120812
transform 1 0 1784 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_390
timestamp 1543120812
transform 1 0 1704 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_391
timestamp 1543120812
transform 1 0 2296 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_392
timestamp 1543120812
transform 1 0 2216 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_393
timestamp 1543120812
transform 1 0 1560 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_394
timestamp 1543120812
transform 1 0 1480 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_395
timestamp 1543120812
transform 1 0 808 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_396
timestamp 1543120812
transform 1 0 744 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_397
timestamp 1543120812
transform 1 0 2104 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_398
timestamp 1543120812
transform 1 0 2024 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_399
timestamp 1543120812
transform 1 0 2136 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_400
timestamp 1543120812
transform 1 0 2008 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_401
timestamp 1543120812
transform 1 0 1336 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_402
timestamp 1543120812
transform 1 0 1288 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_403
timestamp 1543120812
transform 1 0 1640 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_404
timestamp 1543120812
transform 1 0 1576 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_405
timestamp 1543120812
transform 1 0 2360 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_406
timestamp 1543120812
transform 1 0 2088 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_407
timestamp 1543120812
transform 1 0 3128 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_408
timestamp 1543120812
transform 1 0 2968 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_409
timestamp 1543120812
transform 1 0 2648 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_410
timestamp 1543120812
transform 1 0 2120 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_411
timestamp 1543120812
transform 1 0 2104 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_412
timestamp 1543120812
transform 1 0 1992 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_413
timestamp 1543120812
transform 1 0 1624 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_414
timestamp 1543120812
transform 1 0 1511 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_415
timestamp 1543120812
transform 1 0 1240 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_416
timestamp 1543120812
transform 1 0 888 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_417
timestamp 1543120812
transform 1 0 616 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_418
timestamp 1543120812
transform 1 0 1560 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_419
timestamp 1543120812
transform 1 0 1320 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_420
timestamp 1543120812
transform 1 0 1160 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_421
timestamp 1543120812
transform 1 0 984 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_422
timestamp 1543120812
transform 1 0 696 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_423
timestamp 1543120812
transform 1 0 3352 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_424
timestamp 1543120812
transform 1 0 3224 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_425
timestamp 1543120812
transform 1 0 2792 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_426
timestamp 1543120812
transform 1 0 2376 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_427
timestamp 1543120812
transform 1 0 2264 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_428
timestamp 1543120812
transform 1 0 2248 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_429
timestamp 1543120812
transform 1 0 584 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_430
timestamp 1543120812
transform 1 0 552 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_431
timestamp 1543120812
transform 1 0 424 0 1 3010
box -4 -4 4 4
use M2_M1  M2_M1_432
timestamp 1543120812
transform 1 0 424 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_433
timestamp 1543120812
transform 1 0 2248 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_434
timestamp 1543120812
transform 1 0 2136 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_435
timestamp 1543120812
transform 1 0 2632 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_436
timestamp 1543120812
transform 1 0 2504 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_437
timestamp 1543120812
transform 1 0 680 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_438
timestamp 1543120812
transform 1 0 552 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_439
timestamp 1543120812
transform 1 0 3160 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_440
timestamp 1543120812
transform 1 0 2952 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_441
timestamp 1543120812
transform 1 0 2648 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_442
timestamp 1543120812
transform 1 0 2424 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_443
timestamp 1543120812
transform 1 0 2376 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_444
timestamp 1543120812
transform 1 0 1048 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_445
timestamp 1543120812
transform 1 0 968 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_446
timestamp 1543120812
transform 1 0 776 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_447
timestamp 1543120812
transform 1 0 776 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_448
timestamp 1543120812
transform 1 0 1272 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_449
timestamp 1543120812
transform 1 0 1080 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_450
timestamp 1543120812
transform 1 0 1080 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_451
timestamp 1543120812
transform 1 0 1048 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_452
timestamp 1543120812
transform 1 0 3016 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_453
timestamp 1543120812
transform 1 0 2536 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_454
timestamp 1543120812
transform 1 0 2536 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_455
timestamp 1543120812
transform 1 0 2520 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_456
timestamp 1543120812
transform 1 0 1016 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_457
timestamp 1543120812
transform 1 0 968 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_458
timestamp 1543120812
transform 1 0 2872 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_459
timestamp 1543120812
transform 1 0 2632 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_460
timestamp 1543120812
transform 1 0 2392 0 1 2390
box -4 -4 4 4
use M2_M1  M2_M1_461
timestamp 1543120812
transform 1 0 2376 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_462
timestamp 1543120812
transform 1 0 2376 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_463
timestamp 1543120812
transform 1 0 1784 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_464
timestamp 1543120812
transform 1 0 1752 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_465
timestamp 1543120812
transform 1 0 1256 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_466
timestamp 1543120812
transform 1 0 808 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_467
timestamp 1543120812
transform 1 0 696 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_468
timestamp 1543120812
transform 1 0 1672 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_469
timestamp 1543120812
transform 1 0 1640 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_470
timestamp 1543120812
transform 1 0 1432 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_471
timestamp 1543120812
transform 1 0 1208 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_472
timestamp 1543120812
transform 1 0 888 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_473
timestamp 1543120812
transform 1 0 3272 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_474
timestamp 1543120812
transform 1 0 2968 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_475
timestamp 1543120812
transform 1 0 2760 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_476
timestamp 1543120812
transform 1 0 2552 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_477
timestamp 1543120812
transform 1 0 2536 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_478
timestamp 1543120812
transform 1 0 2520 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_479
timestamp 1543120812
transform 1 0 1752 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_480
timestamp 1543120812
transform 1 0 1640 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_481
timestamp 1543120812
transform 1 0 1608 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_482
timestamp 1543120812
transform 1 0 1000 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_483
timestamp 1543120812
transform 1 0 872 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_484
timestamp 1543120812
transform 1 0 1688 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_485
timestamp 1543120812
transform 1 0 1640 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_486
timestamp 1543120812
transform 1 0 1592 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_487
timestamp 1543120812
transform 1 0 1592 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_488
timestamp 1543120812
transform 1 0 1560 0 1 290
box -4 -4 4 4
use M2_M1  M2_M1_489
timestamp 1543120812
transform 1 0 1512 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_490
timestamp 1543120812
transform 1 0 1512 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_491
timestamp 1543120812
transform 1 0 2872 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_492
timestamp 1543120812
transform 1 0 2824 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_493
timestamp 1543120812
transform 1 0 2600 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_494
timestamp 1543120812
transform 1 0 2600 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_495
timestamp 1543120812
transform 1 0 2424 0 1 770
box -4 -4 4 4
use M2_M1  M2_M1_496
timestamp 1543120812
transform 1 0 2088 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_497
timestamp 1543120812
transform 1 0 1816 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_498
timestamp 1543120812
transform 1 0 1448 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_499
timestamp 1543120812
transform 1 0 1416 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_500
timestamp 1543120812
transform 1 0 1304 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_501
timestamp 1543120812
transform 1 0 1112 0 1 1650
box -4 -4 4 4
use M2_M1  M2_M1_502
timestamp 1543120812
transform 1 0 1112 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_503
timestamp 1543120812
transform 1 0 872 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_504
timestamp 1543120812
transform 1 0 632 0 1 1830
box -4 -4 4 4
use M2_M1  M2_M1_505
timestamp 1543120812
transform 1 0 600 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_506
timestamp 1543120812
transform 1 0 984 0 1 790
box -4 -4 4 4
use M2_M1  M2_M1_507
timestamp 1543120812
transform 1 0 920 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_508
timestamp 1543120812
transform 1 0 2536 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_509
timestamp 1543120812
transform 1 0 2488 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_510
timestamp 1543120812
transform 1 0 2360 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_511
timestamp 1543120812
transform 1 0 1784 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_512
timestamp 1543120812
transform 1 0 1784 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_513
timestamp 1543120812
transform 1 0 2280 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_514
timestamp 1543120812
transform 1 0 2280 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_515
timestamp 1543120812
transform 1 0 1896 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_516
timestamp 1543120812
transform 1 0 1768 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_517
timestamp 1543120812
transform 1 0 1768 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_518
timestamp 1543120812
transform 1 0 1320 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_519
timestamp 1543120812
transform 1 0 1320 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_520
timestamp 1543120812
transform 1 0 2280 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_521
timestamp 1543120812
transform 1 0 2088 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_522
timestamp 1543120812
transform 1 0 1992 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_523
timestamp 1543120812
transform 1 0 1544 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_524
timestamp 1543120812
transform 1 0 1272 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_525
timestamp 1543120812
transform 1 0 2136 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_526
timestamp 1543120812
transform 1 0 2056 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_527
timestamp 1543120812
transform 1 0 1800 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_528
timestamp 1543120812
transform 1 0 1624 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_529
timestamp 1543120812
transform 1 0 1432 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_530
timestamp 1543120812
transform 1 0 696 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_531
timestamp 1543120812
transform 1 0 648 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_532
timestamp 1543120812
transform 1 0 2152 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_533
timestamp 1543120812
transform 1 0 2104 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_534
timestamp 1543120812
transform 1 0 1656 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_535
timestamp 1543120812
transform 1 0 1656 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_536
timestamp 1543120812
transform 1 0 1608 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_537
timestamp 1543120812
transform 1 0 1144 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_538
timestamp 1543120812
transform 1 0 1048 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_539
timestamp 1543120812
transform 1 0 904 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_540
timestamp 1543120812
transform 1 0 728 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_541
timestamp 1543120812
transform 1 0 728 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_542
timestamp 1543120812
transform 1 0 1176 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_543
timestamp 1543120812
transform 1 0 1144 0 1 610
box -4 -4 4 4
use M2_M1  M2_M1_544
timestamp 1543120812
transform 1 0 792 0 1 610
box -4 -4 4 4
use M2_M1  M2_M1_545
timestamp 1543120812
transform 1 0 776 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_546
timestamp 1543120812
transform 1 0 456 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_547
timestamp 1543120812
transform 1 0 2728 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_548
timestamp 1543120812
transform 1 0 2648 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_549
timestamp 1543120812
transform 1 0 2040 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_550
timestamp 1543120812
transform 1 0 1960 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_551
timestamp 1543120812
transform 1 0 1992 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_552
timestamp 1543120812
transform 1 0 1992 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_553
timestamp 1543120812
transform 1 0 2360 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_554
timestamp 1543120812
transform 1 0 2280 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_555
timestamp 1543120812
transform 1 0 3336 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_556
timestamp 1543120812
transform 1 0 3304 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_557
timestamp 1543120812
transform 1 0 728 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_558
timestamp 1543120812
transform 1 0 680 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_559
timestamp 1543120812
transform 1 0 648 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_560
timestamp 1543120812
transform 1 0 584 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_561
timestamp 1543120812
transform 1 0 3080 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_562
timestamp 1543120812
transform 1 0 3048 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_563
timestamp 1543120812
transform 1 0 3000 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_564
timestamp 1543120812
transform 1 0 2952 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_565
timestamp 1543120812
transform 1 0 920 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_566
timestamp 1543120812
transform 1 0 872 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_567
timestamp 1543120812
transform 1 0 728 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_568
timestamp 1543120812
transform 1 0 680 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_569
timestamp 1543120812
transform 1 0 3016 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_570
timestamp 1543120812
transform 1 0 2984 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_571
timestamp 1543120812
transform 1 0 3112 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_572
timestamp 1543120812
transform 1 0 3080 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_573
timestamp 1543120812
transform 1 0 1224 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_574
timestamp 1543120812
transform 1 0 1192 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_575
timestamp 1543120812
transform 1 0 808 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_576
timestamp 1543120812
transform 1 0 728 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_577
timestamp 1543120812
transform 1 0 3256 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_578
timestamp 1543120812
transform 1 0 3224 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_579
timestamp 1543120812
transform 1 0 2536 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_580
timestamp 1543120812
transform 1 0 2472 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_581
timestamp 1543120812
transform 1 0 3160 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_582
timestamp 1543120812
transform 1 0 3128 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_583
timestamp 1543120812
transform 1 0 2872 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_584
timestamp 1543120812
transform 1 0 2840 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_585
timestamp 1543120812
transform 1 0 2200 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_586
timestamp 1543120812
transform 1 0 2168 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_587
timestamp 1543120812
transform 1 0 1752 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_588
timestamp 1543120812
transform 1 0 1480 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_589
timestamp 1543120812
transform 1 0 1336 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_590
timestamp 1543120812
transform 1 0 1256 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_591
timestamp 1543120812
transform 1 0 2296 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_592
timestamp 1543120812
transform 1 0 2264 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_593
timestamp 1543120812
transform 1 0 2616 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_594
timestamp 1543120812
transform 1 0 2584 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_595
timestamp 1543120812
transform 1 0 2360 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_596
timestamp 1543120812
transform 1 0 2280 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_597
timestamp 1543120812
transform 1 0 2264 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_598
timestamp 1543120812
transform 1 0 1816 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_599
timestamp 1543120812
transform 1 0 1800 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_600
timestamp 1543120812
transform 1 0 1688 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_601
timestamp 1543120812
transform 1 0 1464 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_602
timestamp 1543120812
transform 1 0 1304 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_603
timestamp 1543120812
transform 1 0 1176 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_604
timestamp 1543120812
transform 1 0 1160 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_605
timestamp 1543120812
transform 1 0 680 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_606
timestamp 1543120812
transform 1 0 344 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_607
timestamp 1543120812
transform 1 0 344 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_608
timestamp 1543120812
transform 1 0 3064 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_609
timestamp 1543120812
transform 1 0 3016 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_610
timestamp 1543120812
transform 1 0 2984 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_611
timestamp 1543120812
transform 1 0 2968 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_612
timestamp 1543120812
transform 1 0 2968 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_613
timestamp 1543120812
transform 1 0 2856 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_614
timestamp 1543120812
transform 1 0 2776 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_615
timestamp 1543120812
transform 1 0 2728 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_616
timestamp 1543120812
transform 1 0 2552 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_617
timestamp 1543120812
transform 1 0 2360 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_618
timestamp 1543120812
transform 1 0 2344 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_619
timestamp 1543120812
transform 1 0 2184 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_620
timestamp 1543120812
transform 1 0 1896 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_621
timestamp 1543120812
transform 1 0 1864 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_622
timestamp 1543120812
transform 1 0 1672 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_623
timestamp 1543120812
transform 1 0 3320 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_624
timestamp 1543120812
transform 1 0 3240 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_625
timestamp 1543120812
transform 1 0 3144 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_626
timestamp 1543120812
transform 1 0 3096 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_627
timestamp 1543120812
transform 1 0 3064 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_628
timestamp 1543120812
transform 1 0 3032 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_629
timestamp 1543120812
transform 1 0 3000 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_630
timestamp 1543120812
transform 1 0 2856 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_631
timestamp 1543120812
transform 1 0 2840 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_632
timestamp 1543120812
transform 1 0 2552 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_633
timestamp 1543120812
transform 1 0 2184 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_634
timestamp 1543120812
transform 1 0 1208 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_635
timestamp 1543120812
transform 1 0 936 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_636
timestamp 1543120812
transform 1 0 920 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_637
timestamp 1543120812
transform 1 0 824 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_638
timestamp 1543120812
transform 1 0 744 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_639
timestamp 1543120812
transform 1 0 744 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_640
timestamp 1543120812
transform 1 0 664 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_641
timestamp 1543120812
transform 1 0 968 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_642
timestamp 1543120812
transform 1 0 936 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_643
timestamp 1543120812
transform 1 0 3176 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_644
timestamp 1543120812
transform 1 0 3160 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_645
timestamp 1543120812
transform 1 0 3080 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_646
timestamp 1543120812
transform 1 0 3032 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_647
timestamp 1543120812
transform 1 0 3000 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_648
timestamp 1543120812
transform 1 0 2952 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_649
timestamp 1543120812
transform 1 0 2952 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_650
timestamp 1543120812
transform 1 0 2920 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_651
timestamp 1543120812
transform 1 0 2920 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_652
timestamp 1543120812
transform 1 0 2744 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_653
timestamp 1543120812
transform 1 0 2488 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_654
timestamp 1543120812
transform 1 0 1976 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_655
timestamp 1543120812
transform 1 0 1144 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_656
timestamp 1543120812
transform 1 0 872 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_657
timestamp 1543120812
transform 1 0 760 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_658
timestamp 1543120812
transform 1 0 760 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_659
timestamp 1543120812
transform 1 0 680 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_660
timestamp 1543120812
transform 1 0 616 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_661
timestamp 1543120812
transform 1 0 600 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_662
timestamp 1543120812
transform 1 0 3160 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_663
timestamp 1543120812
transform 1 0 3080 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_664
timestamp 1543120812
transform 1 0 3080 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_665
timestamp 1543120812
transform 1 0 3000 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_666
timestamp 1543120812
transform 1 0 2984 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_667
timestamp 1543120812
transform 1 0 2936 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_668
timestamp 1543120812
transform 1 0 2824 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_669
timestamp 1543120812
transform 1 0 2776 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_670
timestamp 1543120812
transform 1 0 2680 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_671
timestamp 1543120812
transform 1 0 2440 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_672
timestamp 1543120812
transform 1 0 2056 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_673
timestamp 1543120812
transform 1 0 1640 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_674
timestamp 1543120812
transform 1 0 1448 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_675
timestamp 1543120812
transform 1 0 1080 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_676
timestamp 1543120812
transform 1 0 968 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_677
timestamp 1543120812
transform 1 0 856 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_678
timestamp 1543120812
transform 1 0 808 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_679
timestamp 1543120812
transform 1 0 696 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_680
timestamp 1543120812
transform 1 0 616 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_681
timestamp 1543120812
transform 1 0 3240 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_682
timestamp 1543120812
transform 1 0 3208 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_683
timestamp 1543120812
transform 1 0 2440 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_684
timestamp 1543120812
transform 1 0 2376 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_685
timestamp 1543120812
transform 1 0 2712 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_686
timestamp 1543120812
transform 1 0 2648 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_687
timestamp 1543120812
transform 1 0 2792 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_688
timestamp 1543120812
transform 1 0 2728 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_689
timestamp 1543120812
transform 1 0 2984 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_690
timestamp 1543120812
transform 1 0 2920 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_691
timestamp 1543120812
transform 1 0 3592 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_692
timestamp 1543120812
transform 1 0 3528 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_693
timestamp 1543120812
transform 1 0 3416 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_694
timestamp 1543120812
transform 1 0 3352 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_695
timestamp 1543120812
transform 1 0 3608 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_696
timestamp 1543120812
transform 1 0 3608 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_697
timestamp 1543120812
transform 1 0 3640 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_698
timestamp 1543120812
transform 1 0 3576 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_699
timestamp 1543120812
transform 1 0 3480 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_700
timestamp 1543120812
transform 1 0 3368 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_701
timestamp 1543120812
transform 1 0 3480 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_702
timestamp 1543120812
transform 1 0 3368 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_703
timestamp 1543120812
transform 1 0 2856 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_704
timestamp 1543120812
transform 1 0 2856 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_705
timestamp 1543120812
transform 1 0 2952 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_706
timestamp 1543120812
transform 1 0 2824 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_707
timestamp 1543120812
transform 1 0 3016 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_708
timestamp 1543120812
transform 1 0 2936 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_709
timestamp 1543120812
transform 1 0 3208 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_710
timestamp 1543120812
transform 1 0 3080 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_711
timestamp 1543120812
transform 1 0 3192 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_712
timestamp 1543120812
transform 1 0 3064 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_713
timestamp 1543120812
transform 1 0 3160 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_714
timestamp 1543120812
transform 1 0 3160 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_715
timestamp 1543120812
transform 1 0 3080 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_716
timestamp 1543120812
transform 1 0 2952 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_717
timestamp 1543120812
transform 1 0 3144 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_718
timestamp 1543120812
transform 1 0 3112 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_719
timestamp 1543120812
transform 1 0 2472 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_720
timestamp 1543120812
transform 1 0 2360 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_721
timestamp 1543120812
transform 1 0 2120 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_722
timestamp 1543120812
transform 1 0 2056 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_723
timestamp 1543120812
transform 1 0 2040 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_724
timestamp 1543120812
transform 1 0 1928 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_725
timestamp 1543120812
transform 1 0 2728 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_726
timestamp 1543120812
transform 1 0 2616 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_727
timestamp 1543120812
transform 1 0 2936 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_728
timestamp 1543120812
transform 1 0 2840 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_729
timestamp 1543120812
transform 1 0 3064 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_730
timestamp 1543120812
transform 1 0 2888 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_731
timestamp 1543120812
transform 1 0 2984 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_732
timestamp 1543120812
transform 1 0 2984 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_733
timestamp 1543120812
transform 1 0 1944 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_734
timestamp 1543120812
transform 1 0 1912 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_735
timestamp 1543120812
transform 1 0 1736 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_736
timestamp 1543120812
transform 1 0 2024 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_737
timestamp 1543120812
transform 1 0 1928 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_738
timestamp 1543120812
transform 1 0 1848 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_739
timestamp 1543120812
transform 1 0 2024 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_740
timestamp 1543120812
transform 1 0 1864 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_741
timestamp 1543120812
transform 1 0 1864 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_742
timestamp 1543120812
transform 1 0 1944 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_743
timestamp 1543120812
transform 1 0 1800 0 1 3430
box -4 -4 4 4
use M2_M1  M2_M1_744
timestamp 1543120812
transform 1 0 1800 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_745
timestamp 1543120812
transform 1 0 1608 0 1 3430
box -4 -4 4 4
use M2_M1  M2_M1_746
timestamp 1543120812
transform 1 0 1800 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_747
timestamp 1543120812
transform 1 0 1784 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_748
timestamp 1543120812
transform 1 0 1768 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_749
timestamp 1543120812
transform 1 0 1624 0 1 3410
box -4 -4 4 4
use M2_M1  M2_M1_750
timestamp 1543120812
transform 1 0 792 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_751
timestamp 1543120812
transform 1 0 568 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_752
timestamp 1543120812
transform 1 0 424 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_753
timestamp 1543120812
transform 1 0 648 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_754
timestamp 1543120812
transform 1 0 616 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_755
timestamp 1543120812
transform 1 0 616 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_756
timestamp 1543120812
transform 1 0 408 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_757
timestamp 1543120812
transform 1 0 2072 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_758
timestamp 1543120812
transform 1 0 1928 0 1 1990
box -4 -4 4 4
use M2_M1  M2_M1_759
timestamp 1543120812
transform 1 0 1928 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_760
timestamp 1543120812
transform 1 0 1560 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_761
timestamp 1543120812
transform 1 0 1240 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_762
timestamp 1543120812
transform 1 0 1128 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_763
timestamp 1543120812
transform 1 0 1768 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_764
timestamp 1543120812
transform 1 0 1752 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_765
timestamp 1543120812
transform 1 0 1608 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_766
timestamp 1543120812
transform 1 0 1592 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_767
timestamp 1543120812
transform 1 0 1528 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_768
timestamp 1543120812
transform 1 0 1768 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_769
timestamp 1543120812
transform 1 0 1752 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_770
timestamp 1543120812
transform 1 0 1640 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_771
timestamp 1543120812
transform 1 0 1336 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_772
timestamp 1543120812
transform 1 0 1240 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_773
timestamp 1543120812
transform 1 0 2472 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_774
timestamp 1543120812
transform 1 0 2264 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_775
timestamp 1543120812
transform 1 0 2152 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_776
timestamp 1543120812
transform 1 0 2072 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_777
timestamp 1543120812
transform 1 0 2040 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_778
timestamp 1543120812
transform 1 0 2184 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_779
timestamp 1543120812
transform 1 0 2040 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_780
timestamp 1543120812
transform 1 0 1992 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_781
timestamp 1543120812
transform 1 0 1496 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_782
timestamp 1543120812
transform 1 0 1304 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_783
timestamp 1543120812
transform 1 0 1208 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_784
timestamp 1543120812
transform 1 0 2520 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_785
timestamp 1543120812
transform 1 0 2264 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_786
timestamp 1543120812
transform 1 0 2264 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_787
timestamp 1543120812
transform 1 0 2216 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_788
timestamp 1543120812
transform 1 0 2120 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_789
timestamp 1543120812
transform 1 0 1304 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_790
timestamp 1543120812
transform 1 0 1256 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_791
timestamp 1543120812
transform 1 0 1496 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_792
timestamp 1543120812
transform 1 0 1352 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_793
timestamp 1543120812
transform 1 0 1256 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_794
timestamp 1543120812
transform 1 0 1160 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_795
timestamp 1543120812
transform 1 0 1336 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_796
timestamp 1543120812
transform 1 0 1288 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_797
timestamp 1543120812
transform 1 0 1240 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_798
timestamp 1543120812
transform 1 0 2232 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_799
timestamp 1543120812
transform 1 0 2232 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_800
timestamp 1543120812
transform 1 0 1928 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_801
timestamp 1543120812
transform 1 0 1720 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_802
timestamp 1543120812
transform 1 0 1720 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_803
timestamp 1543120812
transform 1 0 1608 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_804
timestamp 1543120812
transform 1 0 1560 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_805
timestamp 1543120812
transform 1 0 2472 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_806
timestamp 1543120812
transform 1 0 2392 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_807
timestamp 1543120812
transform 1 0 2392 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_808
timestamp 1543120812
transform 1 0 1736 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_809
timestamp 1543120812
transform 1 0 1736 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_810
timestamp 1543120812
transform 1 0 1192 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_811
timestamp 1543120812
transform 1 0 1000 0 1 870
box -4 -4 4 4
use M2_M1  M2_M1_812
timestamp 1543120812
transform 1 0 984 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_813
timestamp 1543120812
transform 1 0 984 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_814
timestamp 1543120812
transform 1 0 856 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_815
timestamp 1543120812
transform 1 0 824 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_816
timestamp 1543120812
transform 1 0 952 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_817
timestamp 1543120812
transform 1 0 936 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_818
timestamp 1543120812
transform 1 0 936 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_819
timestamp 1543120812
transform 1 0 904 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_820
timestamp 1543120812
transform 1 0 888 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_821
timestamp 1543120812
transform 1 0 696 0 1 1650
box -4 -4 4 4
use M2_M1  M2_M1_822
timestamp 1543120812
transform 1 0 648 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_823
timestamp 1543120812
transform 1 0 872 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_824
timestamp 1543120812
transform 1 0 760 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_825
timestamp 1543120812
transform 1 0 632 0 1 1650
box -4 -4 4 4
use M2_M1  M2_M1_826
timestamp 1543120812
transform 1 0 568 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_827
timestamp 1543120812
transform 1 0 904 0 1 1650
box -4 -4 4 4
use M2_M1  M2_M1_828
timestamp 1543120812
transform 1 0 600 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_829
timestamp 1543120812
transform 1 0 600 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_830
timestamp 1543120812
transform 1 0 760 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_831
timestamp 1543120812
transform 1 0 600 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_832
timestamp 1543120812
transform 1 0 520 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_833
timestamp 1543120812
transform 1 0 520 0 1 690
box -4 -4 4 4
use M2_M1  M2_M1_834
timestamp 1543120812
transform 1 0 568 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_835
timestamp 1543120812
transform 1 0 504 0 1 850
box -4 -4 4 4
use M2_M1  M2_M1_836
timestamp 1543120812
transform 1 0 808 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_837
timestamp 1543120812
transform 1 0 808 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_838
timestamp 1543120812
transform 1 0 472 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_839
timestamp 1543120812
transform 1 0 520 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_840
timestamp 1543120812
transform 1 0 488 0 1 870
box -4 -4 4 4
use M2_M1  M2_M1_841
timestamp 1543120812
transform 1 0 1224 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_842
timestamp 1543120812
transform 1 0 1160 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_843
timestamp 1543120812
transform 1 0 936 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_844
timestamp 1543120812
transform 1 0 728 0 1 630
box -4 -4 4 4
use M2_M1  M2_M1_845
timestamp 1543120812
transform 1 0 792 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_846
timestamp 1543120812
transform 1 0 760 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_847
timestamp 1543120812
transform 1 0 1016 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_848
timestamp 1543120812
transform 1 0 744 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_849
timestamp 1543120812
transform 1 0 824 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_850
timestamp 1543120812
transform 1 0 728 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_851
timestamp 1543120812
transform 1 0 696 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_852
timestamp 1543120812
transform 1 0 680 0 1 1190
box -4 -4 4 4
use M2_M1  M2_M1_853
timestamp 1543120812
transform 1 0 792 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_854
timestamp 1543120812
transform 1 0 792 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_855
timestamp 1543120812
transform 1 0 1368 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_856
timestamp 1543120812
transform 1 0 1176 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_857
timestamp 1543120812
transform 1 0 968 0 1 1090
box -4 -4 4 4
use M2_M1  M2_M1_858
timestamp 1543120812
transform 1 0 840 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_859
timestamp 1543120812
transform 1 0 840 0 1 1090
box -4 -4 4 4
use M2_M1  M2_M1_860
timestamp 1543120812
transform 1 0 824 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_861
timestamp 1543120812
transform 1 0 792 0 1 1490
box -4 -4 4 4
use M2_M1  M2_M1_862
timestamp 1543120812
transform 1 0 632 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_863
timestamp 1543120812
transform 1 0 632 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_864
timestamp 1543120812
transform 1 0 616 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_865
timestamp 1543120812
transform 1 0 1288 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_866
timestamp 1543120812
transform 1 0 968 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_867
timestamp 1543120812
transform 1 0 792 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_868
timestamp 1543120812
transform 1 0 1192 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_869
timestamp 1543120812
transform 1 0 952 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_870
timestamp 1543120812
transform 1 0 1800 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_871
timestamp 1543120812
transform 1 0 1208 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_872
timestamp 1543120812
transform 1 0 1208 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_873
timestamp 1543120812
transform 1 0 1112 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_874
timestamp 1543120812
transform 1 0 1080 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_875
timestamp 1543120812
transform 1 0 1112 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_876
timestamp 1543120812
transform 1 0 1112 0 1 870
box -4 -4 4 4
use M2_M1  M2_M1_877
timestamp 1543120812
transform 1 0 1000 0 1 1250
box -4 -4 4 4
use M2_M1  M2_M1_878
timestamp 1543120812
transform 1 0 968 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_879
timestamp 1543120812
transform 1 0 1016 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_880
timestamp 1543120812
transform 1 0 968 0 1 1270
box -4 -4 4 4
use M2_M1  M2_M1_881
timestamp 1543120812
transform 1 0 1928 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_882
timestamp 1543120812
transform 1 0 1240 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_883
timestamp 1543120812
transform 1 0 1416 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_884
timestamp 1543120812
transform 1 0 1256 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_885
timestamp 1543120812
transform 1 0 1288 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_886
timestamp 1543120812
transform 1 0 1288 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_887
timestamp 1543120812
transform 1 0 1496 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_888
timestamp 1543120812
transform 1 0 1416 0 1 1030
box -4 -4 4 4
use M2_M1  M2_M1_889
timestamp 1543120812
transform 1 0 1576 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_890
timestamp 1543120812
transform 1 0 1464 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_891
timestamp 1543120812
transform 1 0 1960 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_892
timestamp 1543120812
transform 1 0 1480 0 1 1010
box -4 -4 4 4
use M2_M1  M2_M1_893
timestamp 1543120812
transform 1 0 2104 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_894
timestamp 1543120812
transform 1 0 1992 0 1 1090
box -4 -4 4 4
use M2_M1  M2_M1_895
timestamp 1543120812
transform 1 0 2056 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_896
timestamp 1543120812
transform 1 0 2024 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_897
timestamp 1543120812
transform 1 0 1880 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_898
timestamp 1543120812
transform 1 0 1768 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_899
timestamp 1543120812
transform 1 0 2568 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_900
timestamp 1543120812
transform 1 0 1784 0 1 1410
box -4 -4 4 4
use M2_M1  M2_M1_901
timestamp 1543120812
transform 1 0 2664 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_902
timestamp 1543120812
transform 1 0 2600 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_903
timestamp 1543120812
transform 1 0 1544 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_904
timestamp 1543120812
transform 1 0 1432 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_905
timestamp 1543120812
transform 1 0 1464 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_906
timestamp 1543120812
transform 1 0 1384 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_907
timestamp 1543120812
transform 1 0 2200 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_908
timestamp 1543120812
transform 1 0 1976 0 1 1470
box -4 -4 4 4
use M2_M1  M2_M1_909
timestamp 1543120812
transform 1 0 2088 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_910
timestamp 1543120812
transform 1 0 2008 0 1 1430
box -4 -4 4 4
use M2_M1  M2_M1_911
timestamp 1543120812
transform 1 0 456 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_912
timestamp 1543120812
transform 1 0 360 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_913
timestamp 1543120812
transform 1 0 1640 0 1 3430
box -4 -4 4 4
use M2_M1  M2_M1_914
timestamp 1543120812
transform 1 0 1480 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_915
timestamp 1543120812
transform 1 0 1752 0 1 3450
box -4 -4 4 4
use M2_M1  M2_M1_916
timestamp 1543120812
transform 1 0 1656 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_917
timestamp 1543120812
transform 1 0 1880 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_918
timestamp 1543120812
transform 1 0 1704 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_919
timestamp 1543120812
transform 1 0 1976 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_920
timestamp 1543120812
transform 1 0 1896 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_921
timestamp 1543120812
transform 1 0 1848 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_922
timestamp 1543120812
transform 1 0 2168 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_923
timestamp 1543120812
transform 1 0 1736 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_924
timestamp 1543120812
transform 1 0 1784 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_925
timestamp 1543120812
transform 1 0 1768 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_926
timestamp 1543120812
transform 1 0 1736 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_927
timestamp 1543120812
transform 1 0 1624 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_928
timestamp 1543120812
transform 1 0 2536 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_929
timestamp 1543120812
transform 1 0 1752 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_930
timestamp 1543120812
transform 1 0 1800 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_931
timestamp 1543120812
transform 1 0 1224 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_932
timestamp 1543120812
transform 1 0 2776 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_933
timestamp 1543120812
transform 1 0 1816 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_934
timestamp 1543120812
transform 1 0 2792 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_935
timestamp 1543120812
transform 1 0 2648 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_936
timestamp 1543120812
transform 1 0 1192 0 1 2790
box -4 -4 4 4
use M2_M1  M2_M1_937
timestamp 1543120812
transform 1 0 1032 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_938
timestamp 1543120812
transform 1 0 1224 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_939
timestamp 1543120812
transform 1 0 1192 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_940
timestamp 1543120812
transform 1 0 2632 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_941
timestamp 1543120812
transform 1 0 2568 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_942
timestamp 1543120812
transform 1 0 1544 0 1 2290
box -4 -4 4 4
use M2_M1  M2_M1_943
timestamp 1543120812
transform 1 0 1416 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_944
timestamp 1543120812
transform 1 0 1576 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_945
timestamp 1543120812
transform 1 0 1544 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_946
timestamp 1543120812
transform 1 0 1672 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_947
timestamp 1543120812
transform 1 0 1368 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_948
timestamp 1543120812
transform 1 0 2264 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_949
timestamp 1543120812
transform 1 0 2152 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_950
timestamp 1543120812
transform 1 0 2184 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_951
timestamp 1543120812
transform 1 0 2152 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_952
timestamp 1543120812
transform 1 0 1864 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_953
timestamp 1543120812
transform 1 0 1816 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_954
timestamp 1543120812
transform 1 0 1816 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_955
timestamp 1543120812
transform 1 0 1528 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_956
timestamp 1543120812
transform 1 0 1880 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_957
timestamp 1543120812
transform 1 0 1864 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_958
timestamp 1543120812
transform 1 0 1816 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_959
timestamp 1543120812
transform 1 0 1368 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_960
timestamp 1543120812
transform 1 0 1896 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_961
timestamp 1543120812
transform 1 0 1848 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_962
timestamp 1543120812
transform 1 0 1928 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_963
timestamp 1543120812
transform 1 0 1224 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_964
timestamp 1543120812
transform 1 0 2504 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_965
timestamp 1543120812
transform 1 0 1880 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_966
timestamp 1543120812
transform 1 0 2488 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_967
timestamp 1543120812
transform 1 0 2488 0 1 2690
box -4 -4 4 4
use M2_M1  M2_M1_968
timestamp 1543120812
transform 1 0 2600 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_969
timestamp 1543120812
transform 1 0 2536 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_970
timestamp 1543120812
transform 1 0 1192 0 1 2690
box -4 -4 4 4
use M2_M1  M2_M1_971
timestamp 1543120812
transform 1 0 920 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_972
timestamp 1543120812
transform 1 0 1224 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_973
timestamp 1543120812
transform 1 0 1192 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_974
timestamp 1543120812
transform 1 0 2056 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_975
timestamp 1543120812
transform 1 0 1944 0 1 2690
box -4 -4 4 4
use M2_M1  M2_M1_976
timestamp 1543120812
transform 1 0 2440 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_977
timestamp 1543120812
transform 1 0 1992 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_978
timestamp 1543120812
transform 1 0 1384 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_979
timestamp 1543120812
transform 1 0 1336 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_980
timestamp 1543120812
transform 1 0 1480 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_981
timestamp 1543120812
transform 1 0 1464 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_982
timestamp 1543120812
transform 1 0 1512 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_983
timestamp 1543120812
transform 1 0 1480 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_984
timestamp 1543120812
transform 1 0 2376 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_985
timestamp 1543120812
transform 1 0 1880 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_986
timestamp 1543120812
transform 1 0 1992 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_987
timestamp 1543120812
transform 1 0 1912 0 1 2850
box -4 -4 4 4
use M2_M1  M2_M1_988
timestamp 1543120812
transform 1 0 2232 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_989
timestamp 1543120812
transform 1 0 1976 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_990
timestamp 1543120812
transform 1 0 1944 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_991
timestamp 1543120812
transform 1 0 1896 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_992
timestamp 1543120812
transform 1 0 2024 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_993
timestamp 1543120812
transform 1 0 2008 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_994
timestamp 1543120812
transform 1 0 1928 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_995
timestamp 1543120812
transform 1 0 1544 0 1 2390
box -4 -4 4 4
use M2_M1  M2_M1_996
timestamp 1543120812
transform 1 0 2248 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_997
timestamp 1543120812
transform 1 0 1992 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_998
timestamp 1543120812
transform 1 0 2040 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_999
timestamp 1543120812
transform 1 0 1960 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1000
timestamp 1543120812
transform 1 0 2168 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_1001
timestamp 1543120812
transform 1 0 2104 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1002
timestamp 1543120812
transform 1 0 2440 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1003
timestamp 1543120812
transform 1 0 2328 0 1 2290
box -4 -4 4 4
use M2_M1  M2_M1_1004
timestamp 1543120812
transform 1 0 2584 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1005
timestamp 1543120812
transform 1 0 2360 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1006
timestamp 1543120812
transform 1 0 1928 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1007
timestamp 1543120812
transform 1 0 1784 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1008
timestamp 1543120812
transform 1 0 2344 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1009
timestamp 1543120812
transform 1 0 2280 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1010
timestamp 1543120812
transform 1 0 1576 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1011
timestamp 1543120812
transform 1 0 1448 0 1 2390
box -4 -4 4 4
use M2_M1  M2_M1_1012
timestamp 1543120812
transform 1 0 1480 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1013
timestamp 1543120812
transform 1 0 1448 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1014
timestamp 1543120812
transform 1 0 1880 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1015
timestamp 1543120812
transform 1 0 1736 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1016
timestamp 1543120812
transform 1 0 2328 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1017
timestamp 1543120812
transform 1 0 2216 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1018
timestamp 1543120812
transform 1 0 2248 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1019
timestamp 1543120812
transform 1 0 2216 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1020
timestamp 1543120812
transform 1 0 2648 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1021
timestamp 1543120812
transform 1 0 1896 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1022
timestamp 1543120812
transform 1 0 1912 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1023
timestamp 1543120812
transform 1 0 1592 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1024
timestamp 1543120812
transform 1 0 1944 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1025
timestamp 1543120812
transform 1 0 1864 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1026
timestamp 1543120812
transform 1 0 2776 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_1027
timestamp 1543120812
transform 1 0 1848 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1028
timestamp 1543120812
transform 1 0 1896 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1029
timestamp 1543120812
transform 1 0 1896 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_1030
timestamp 1543120812
transform 1 0 2728 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1031
timestamp 1543120812
transform 1 0 1960 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1032
timestamp 1543120812
transform 1 0 2776 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1033
timestamp 1543120812
transform 1 0 2696 0 1 2390
box -4 -4 4 4
use M2_M1  M2_M1_1034
timestamp 1543120812
transform 1 0 2840 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1035
timestamp 1543120812
transform 1 0 2776 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1036
timestamp 1543120812
transform 1 0 1896 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1037
timestamp 1543120812
transform 1 0 1752 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1038
timestamp 1543120812
transform 1 0 2872 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1039
timestamp 1543120812
transform 1 0 2808 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1040
timestamp 1543120812
transform 1 0 1720 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1041
timestamp 1543120812
transform 1 0 1672 0 1 2390
box -4 -4 4 4
use M2_M1  M2_M1_1042
timestamp 1543120812
transform 1 0 1704 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1043
timestamp 1543120812
transform 1 0 1672 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1044
timestamp 1543120812
transform 1 0 1608 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1045
timestamp 1543120812
transform 1 0 1464 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1046
timestamp 1543120812
transform 1 0 2888 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1047
timestamp 1543120812
transform 1 0 2664 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1048
timestamp 1543120812
transform 1 0 2776 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1049
timestamp 1543120812
transform 1 0 2696 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1050
timestamp 1543120812
transform 1 0 568 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1051
timestamp 1543120812
transform 1 0 472 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1052
timestamp 1543120812
transform 1 0 936 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1053
timestamp 1543120812
transform 1 0 696 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1054
timestamp 1543120812
transform 1 0 648 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1055
timestamp 1543120812
transform 1 0 1528 0 1 3250
box -4 -4 4 4
use M2_M1  M2_M1_1056
timestamp 1543120812
transform 1 0 696 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1057
timestamp 1543120812
transform 1 0 664 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1058
timestamp 1543120812
transform 1 0 1048 0 1 2230
box -4 -4 4 4
use M2_M1  M2_M1_1059
timestamp 1543120812
transform 1 0 984 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1060
timestamp 1543120812
transform 1 0 856 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1061
timestamp 1543120812
transform 1 0 1112 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1062
timestamp 1543120812
transform 1 0 1016 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1063
timestamp 1543120812
transform 1 0 808 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1064
timestamp 1543120812
transform 1 0 1064 0 1 2630
box -4 -4 4 4
use M2_M1  M2_M1_1065
timestamp 1543120812
transform 1 0 552 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_1066
timestamp 1543120812
transform 1 0 520 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_1067
timestamp 1543120812
transform 1 0 1304 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1068
timestamp 1543120812
transform 1 0 1064 0 1 3030
box -4 -4 4 4
use M2_M1  M2_M1_1069
timestamp 1543120812
transform 1 0 1192 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1070
timestamp 1543120812
transform 1 0 1064 0 1 3010
box -4 -4 4 4
use M2_M1  M2_M1_1071
timestamp 1543120812
transform 1 0 2504 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1072
timestamp 1543120812
transform 1 0 1096 0 1 3010
box -4 -4 4 4
use M2_M1  M2_M1_1073
timestamp 1543120812
transform 1 0 2600 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1074
timestamp 1543120812
transform 1 0 2536 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1075
timestamp 1543120812
transform 1 0 1176 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1076
timestamp 1543120812
transform 1 0 1016 0 1 2230
box -4 -4 4 4
use M2_M1  M2_M1_1077
timestamp 1543120812
transform 1 0 2520 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1078
timestamp 1543120812
transform 1 0 1032 0 1 2210
box -4 -4 4 4
use M2_M1  M2_M1_1079
timestamp 1543120812
transform 1 0 2616 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1080
timestamp 1543120812
transform 1 0 2552 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1081
timestamp 1543120812
transform 1 0 1608 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1082
timestamp 1543120812
transform 1 0 1496 0 1 3250
box -4 -4 4 4
use M2_M1  M2_M1_1083
timestamp 1543120812
transform 1 0 2392 0 1 3210
box -4 -4 4 4
use M2_M1  M2_M1_1084
timestamp 1543120812
transform 1 0 1480 0 1 3270
box -4 -4 4 4
use M2_M1  M2_M1_1085
timestamp 1543120812
transform 1 0 2712 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1086
timestamp 1543120812
transform 1 0 2408 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1087
timestamp 1543120812
transform 1 0 1112 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1088
timestamp 1543120812
transform 1 0 1016 0 1 2630
box -4 -4 4 4
use M2_M1  M2_M1_1089
timestamp 1543120812
transform 1 0 2232 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_1090
timestamp 1543120812
transform 1 0 1048 0 1 2610
box -4 -4 4 4
use M2_M1  M2_M1_1091
timestamp 1543120812
transform 1 0 2328 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1092
timestamp 1543120812
transform 1 0 2264 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1093
timestamp 1543120812
transform 1 0 3128 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1094
timestamp 1543120812
transform 1 0 2984 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_1095
timestamp 1543120812
transform 1 0 1016 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1096
timestamp 1543120812
transform 1 0 904 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1097
timestamp 1543120812
transform 1 0 712 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1098
timestamp 1543120812
transform 1 0 664 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1099
timestamp 1543120812
transform 1 0 2968 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1100
timestamp 1543120812
transform 1 0 2776 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1101
timestamp 1543120812
transform 1 0 3064 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_1102
timestamp 1543120812
transform 1 0 2920 0 1 2830
box -4 -4 4 4
use M2_M1  M2_M1_1103
timestamp 1543120812
transform 1 0 1176 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_1104
timestamp 1543120812
transform 1 0 1128 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1105
timestamp 1543120812
transform 1 0 904 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1106
timestamp 1543120812
transform 1 0 792 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1107
timestamp 1543120812
transform 1 0 3208 0 1 3070
box -4 -4 4 4
use M2_M1  M2_M1_1108
timestamp 1543120812
transform 1 0 3080 0 1 3050
box -4 -4 4 4
use M2_M1  M2_M1_1109
timestamp 1543120812
transform 1 0 2520 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_1110
timestamp 1543120812
transform 1 0 2520 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1111
timestamp 1543120812
transform 1 0 3112 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_1112
timestamp 1543120812
transform 1 0 3096 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1113
timestamp 1543120812
transform 1 0 2824 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_1114
timestamp 1543120812
transform 1 0 2824 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1115
timestamp 1543120812
transform 1 0 2152 0 1 3470
box -4 -4 4 4
use M2_M1  M2_M1_1116
timestamp 1543120812
transform 1 0 2152 0 1 3230
box -4 -4 4 4
use M2_M1  M2_M1_1117
timestamp 1543120812
transform 1 0 3288 0 1 2810
box -4 -4 4 4
use M2_M1  M2_M1_1118
timestamp 1543120812
transform 1 0 3256 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1119
timestamp 1543120812
transform 1 0 856 0 1 2430
box -4 -4 4 4
use M2_M1  M2_M1_1120
timestamp 1543120812
transform 1 0 712 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1121
timestamp 1543120812
transform 1 0 744 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1122
timestamp 1543120812
transform 1 0 632 0 1 2670
box -4 -4 4 4
use M2_M1  M2_M1_1123
timestamp 1543120812
transform 1 0 3032 0 1 2650
box -4 -4 4 4
use M2_M1  M2_M1_1124
timestamp 1543120812
transform 1 0 3032 0 1 2410
box -4 -4 4 4
use M2_M1  M2_M1_1125
timestamp 1543120812
transform 1 0 2216 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1126
timestamp 1543120812
transform 1 0 2104 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1127
timestamp 1543120812
transform 1 0 1592 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1128
timestamp 1543120812
transform 1 0 1480 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1129
timestamp 1543120812
transform 1 0 1320 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1130
timestamp 1543120812
transform 1 0 1256 0 1 2030
box -4 -4 4 4
use M2_M1  M2_M1_1131
timestamp 1543120812
transform 1 0 2024 0 1 2250
box -4 -4 4 4
use M2_M1  M2_M1_1132
timestamp 1543120812
transform 1 0 2024 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1133
timestamp 1543120812
transform 1 0 2056 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1134
timestamp 1543120812
transform 1 0 2056 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1135
timestamp 1543120812
transform 1 0 1224 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1136
timestamp 1543120812
transform 1 0 1144 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1137
timestamp 1543120812
transform 1 0 1512 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1138
timestamp 1543120812
transform 1 0 1400 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_1139
timestamp 1543120812
transform 1 0 2312 0 1 1450
box -4 -4 4 4
use M2_M1  M2_M1_1140
timestamp 1543120812
transform 1 0 2248 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1141
timestamp 1543120812
transform 1 0 2424 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_1142
timestamp 1543120812
transform 1 0 2248 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_1143
timestamp 1543120812
transform 1 0 1736 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_1144
timestamp 1543120812
transform 1 0 1736 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_1145
timestamp 1543120812
transform 1 0 1848 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_1146
timestamp 1543120812
transform 1 0 1736 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_1147
timestamp 1543120812
transform 1 0 1752 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1148
timestamp 1543120812
transform 1 0 1560 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1149
timestamp 1543120812
transform 1 0 1864 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_1150
timestamp 1543120812
transform 1 0 1752 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1151
timestamp 1543120812
transform 1 0 2664 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1152
timestamp 1543120812
transform 1 0 2456 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1153
timestamp 1543120812
transform 1 0 2632 0 1 1630
box -4 -4 4 4
use M2_M1  M2_M1_1154
timestamp 1543120812
transform 1 0 2504 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1155
timestamp 1543120812
transform 1 0 728 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1156
timestamp 1543120812
transform 1 0 728 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1157
timestamp 1543120812
transform 1 0 520 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1158
timestamp 1543120812
transform 1 0 440 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_1159
timestamp 1543120812
transform 1 0 568 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_1160
timestamp 1543120812
transform 1 0 440 0 1 1050
box -4 -4 4 4
use M2_M1  M2_M1_1161
timestamp 1543120812
transform 1 0 1240 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1162
timestamp 1543120812
transform 1 0 1240 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_1163
timestamp 1543120812
transform 1 0 744 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_1164
timestamp 1543120812
transform 1 0 744 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_1165
timestamp 1543120812
transform 1 0 2424 0 1 1230
box -4 -4 4 4
use M2_M1  M2_M1_1166
timestamp 1543120812
transform 1 0 2248 0 1 1210
box -4 -4 4 4
use M2_M1  M2_M1_1167
timestamp 1543120812
transform 1 0 1736 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_1168
timestamp 1543120812
transform 1 0 1720 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_1169
timestamp 1543120812
transform 1 0 1528 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_1170
timestamp 1543120812
transform 1 0 1496 0 1 390
box -4 -4 4 4
use M2_M1  M2_M1_1171
timestamp 1543120812
transform 1 0 1480 0 1 230
box -4 -4 4 4
use M2_M1  M2_M1_1172
timestamp 1543120812
transform 1 0 1512 0 1 230
box -4 -4 4 4
use M2_M1  M2_M1_1173
timestamp 1543120812
transform 1 0 1336 0 1 270
box -4 -4 4 4
use M2_M1  M2_M1_1174
timestamp 1543120812
transform 1 0 3176 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_1175
timestamp 1543120812
transform 1 0 3144 0 1 1090
box -4 -4 4 4
use M2_M1  M2_M1_1176
timestamp 1543120812
transform 1 0 3112 0 1 1610
box -4 -4 4 4
use M2_M1  M2_M1_1177
timestamp 1543120812
transform 1 0 3112 0 1 1190
box -4 -4 4 4
use M2_M1  M2_M1_1178
timestamp 1543120812
transform 1 0 3032 0 1 1590
box -4 -4 4 4
use M2_M1  M2_M1_1179
timestamp 1543120812
transform 1 0 2920 0 1 810
box -4 -4 4 4
use M2_M1  M2_M1_1180
timestamp 1543120812
transform 1 0 2856 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1181
timestamp 1543120812
transform 1 0 2632 0 1 1070
box -4 -4 4 4
use M2_M1  M2_M1_1182
timestamp 1543120812
transform 1 0 2520 0 1 830
box -4 -4 4 4
use M2_M1  M2_M1_1183
timestamp 1543120812
transform 1 0 2136 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1184
timestamp 1543120812
transform 1 0 1944 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1185
timestamp 1543120812
transform 1 0 1880 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_1186
timestamp 1543120812
transform 1 0 1080 0 1 1190
box -4 -4 4 4
use M2_M1  M2_M1_1187
timestamp 1543120812
transform 1 0 1608 0 1 650
box -4 -4 4 4
use M2_M1  M2_M1_1188
timestamp 1543120812
transform 1 0 1384 0 1 670
box -4 -4 4 4
use M2_M1  M2_M1_1189
timestamp 1543120812
transform 1 0 1384 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_1190
timestamp 1543120812
transform 1 0 840 0 1 1850
box -4 -4 4 4
use M2_M1  M2_M1_1191
timestamp 1543120812
transform 1 0 600 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1192
timestamp 1543120812
transform 1 0 1832 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_1193
timestamp 1543120812
transform 1 0 1544 0 1 410
box -4 -4 4 4
use M2_M1  M2_M1_1194
timestamp 1543120812
transform 1 0 1448 0 1 430
box -4 -4 4 4
use M2_M1  M2_M1_1195
timestamp 1543120812
transform 1 0 1592 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_1196
timestamp 1543120812
transform 1 0 1320 0 1 250
box -4 -4 4 4
use M2_M1  M2_M1_1197
timestamp 1543120812
transform 1 0 2168 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1198
timestamp 1543120812
transform 1 0 2168 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1199
timestamp 1543120812
transform 1 0 1976 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1200
timestamp 1543120812
transform 1 0 1960 0 1 2270
box -4 -4 4 4
use M2_M1  M2_M1_1201
timestamp 1543120812
transform 1 0 1384 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1202
timestamp 1543120812
transform 1 0 1160 0 1 2010
box -4 -4 4 4
use M2_M1  M2_M1_1203
timestamp 1543120812
transform 1 0 1064 0 1 1870
box -4 -4 4 4
use M2_M1  M2_M1_1204
timestamp 1543120812
transform 1 0 680 0 1 1870
box -4 -4 4 4
use M3_M2  M3_M2_0
timestamp 1543120812
transform 1 0 2744 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_1
timestamp 1543120812
transform 1 0 2552 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_2
timestamp 1543120812
transform 1 0 2280 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_3
timestamp 1543120812
transform 1 0 3160 0 1 330
box -6 -6 6 6
use M3_M2  M3_M2_4
timestamp 1543120812
transform 1 0 2840 0 1 330
box -6 -6 6 6
use M3_M2  M3_M2_5
timestamp 1543120812
transform 1 0 2840 0 1 190
box -6 -6 6 6
use M3_M2  M3_M2_6
timestamp 1543120812
transform 1 0 2632 0 1 190
box -6 -6 6 6
use M3_M2  M3_M2_7
timestamp 1543120812
transform 1 0 3576 0 1 490
box -6 -6 6 6
use M3_M2  M3_M2_8
timestamp 1543120812
transform 1 0 3384 0 1 490
box -6 -6 6 6
use M3_M2  M3_M2_9
timestamp 1543120812
transform 1 0 3256 0 1 490
box -6 -6 6 6
use M3_M2  M3_M2_10
timestamp 1543120812
transform 1 0 3400 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_11
timestamp 1543120812
transform 1 0 3272 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_12
timestamp 1543120812
transform 1 0 3400 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_13
timestamp 1543120812
transform 1 0 3240 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_14
timestamp 1543120812
transform 1 0 2904 0 1 730
box -6 -6 6 6
use M3_M2  M3_M2_15
timestamp 1543120812
transform 1 0 2680 0 1 730
box -6 -6 6 6
use M3_M2  M3_M2_16
timestamp 1543120812
transform 1 0 3288 0 1 890
box -6 -6 6 6
use M3_M2  M3_M2_17
timestamp 1543120812
transform 1 0 3160 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_18
timestamp 1543120812
transform 1 0 3144 0 1 890
box -6 -6 6 6
use M3_M2  M3_M2_19
timestamp 1543120812
transform 1 0 3000 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_20
timestamp 1543120812
transform 1 0 3256 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_21
timestamp 1543120812
transform 1 0 3128 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_22
timestamp 1543120812
transform 1 0 3288 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_23
timestamp 1543120812
transform 1 0 3224 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_24
timestamp 1543120812
transform 1 0 3032 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_25
timestamp 1543120812
transform 1 0 3400 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_26
timestamp 1543120812
transform 1 0 3160 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_27
timestamp 1543120812
transform 1 0 3096 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_28
timestamp 1543120812
transform 1 0 3432 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_29
timestamp 1543120812
transform 1 0 3304 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_30
timestamp 1543120812
transform 1 0 3176 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_31
timestamp 1543120812
transform 1 0 3176 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_32
timestamp 1543120812
transform 1 0 2936 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_33
timestamp 1543120812
transform 1 0 2712 0 1 1290
box -6 -6 6 6
use M3_M2  M3_M2_34
timestamp 1543120812
transform 1 0 2584 0 1 1450
box -6 -6 6 6
use M3_M2  M3_M2_35
timestamp 1543120812
transform 1 0 2584 0 1 1290
box -6 -6 6 6
use M3_M2  M3_M2_36
timestamp 1543120812
transform 1 0 2136 0 1 1450
box -6 -6 6 6
use M3_M2  M3_M2_37
timestamp 1543120812
transform 1 0 2104 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_38
timestamp 1543120812
transform 1 0 1992 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_39
timestamp 1543120812
transform 1 0 1960 0 1 730
box -6 -6 6 6
use M3_M2  M3_M2_40
timestamp 1543120812
transform 1 0 1624 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_41
timestamp 1543120812
transform 1 0 1624 0 1 730
box -6 -6 6 6
use M3_M2  M3_M2_42
timestamp 1543120812
transform 1 0 1544 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_43
timestamp 1543120812
transform 1 0 1432 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_44
timestamp 1543120812
transform 1 0 2136 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_45
timestamp 1543120812
transform 1 0 2056 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_46
timestamp 1543120812
transform 1 0 1816 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_47
timestamp 1543120812
transform 1 0 1512 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_48
timestamp 1543120812
transform 1 0 1464 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_49
timestamp 1543120812
transform 1 0 1448 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_50
timestamp 1543120812
transform 1 0 1320 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_51
timestamp 1543120812
transform 1 0 1320 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_52
timestamp 1543120812
transform 1 0 2504 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_53
timestamp 1543120812
transform 1 0 2440 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_54
timestamp 1543120812
transform 1 0 2424 0 1 810
box -6 -6 6 6
use M3_M2  M3_M2_55
timestamp 1543120812
transform 1 0 2344 0 1 810
box -6 -6 6 6
use M3_M2  M3_M2_56
timestamp 1543120812
transform 1 0 2056 0 1 810
box -6 -6 6 6
use M3_M2  M3_M2_57
timestamp 1543120812
transform 1 0 2024 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_58
timestamp 1543120812
transform 1 0 968 0 1 650
box -6 -6 6 6
use M3_M2  M3_M2_59
timestamp 1543120812
transform 1 0 840 0 1 650
box -6 -6 6 6
use M3_M2  M3_M2_60
timestamp 1543120812
transform 1 0 728 0 1 650
box -6 -6 6 6
use M3_M2  M3_M2_61
timestamp 1543120812
transform 1 0 936 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_62
timestamp 1543120812
transform 1 0 504 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_63
timestamp 1543120812
transform 1 0 1096 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_64
timestamp 1543120812
transform 1 0 1000 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_65
timestamp 1543120812
transform 1 0 1000 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_66
timestamp 1543120812
transform 1 0 680 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_67
timestamp 1543120812
transform 1 0 680 0 1 650
box -6 -6 6 6
use M3_M2  M3_M2_68
timestamp 1543120812
transform 1 0 552 0 1 650
box -6 -6 6 6
use M3_M2  M3_M2_69
timestamp 1543120812
transform 1 0 2920 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_70
timestamp 1543120812
transform 1 0 2904 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_71
timestamp 1543120812
transform 1 0 2760 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_72
timestamp 1543120812
transform 1 0 2680 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_73
timestamp 1543120812
transform 1 0 1960 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_74
timestamp 1543120812
transform 1 0 1960 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_75
timestamp 1543120812
transform 1 0 1784 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_76
timestamp 1543120812
transform 1 0 1784 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_77
timestamp 1543120812
transform 1 0 1736 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_78
timestamp 1543120812
transform 1 0 1688 0 1 1790
box -6 -6 6 6
use M3_M2  M3_M2_79
timestamp 1543120812
transform 1 0 1656 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_80
timestamp 1543120812
transform 1 0 1640 0 1 3130
box -6 -6 6 6
use M3_M2  M3_M2_81
timestamp 1543120812
transform 1 0 1608 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_82
timestamp 1543120812
transform 1 0 1560 0 1 3130
box -6 -6 6 6
use M3_M2  M3_M2_83
timestamp 1543120812
transform 1 0 1560 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_84
timestamp 1543120812
transform 1 0 1512 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_85
timestamp 1543120812
transform 1 0 1512 0 1 1790
box -6 -6 6 6
use M3_M2  M3_M2_86
timestamp 1543120812
transform 1 0 1976 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_87
timestamp 1543120812
transform 1 0 1976 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_88
timestamp 1543120812
transform 1 0 1976 0 1 1510
box -6 -6 6 6
use M3_M2  M3_M2_89
timestamp 1543120812
transform 1 0 1912 0 1 1510
box -6 -6 6 6
use M3_M2  M3_M2_90
timestamp 1543120812
transform 1 0 1896 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_91
timestamp 1543120812
transform 1 0 1848 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_92
timestamp 1543120812
transform 1 0 1848 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_93
timestamp 1543120812
transform 1 0 1752 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_94
timestamp 1543120812
transform 1 0 1736 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_95
timestamp 1543120812
transform 1 0 1688 0 1 1510
box -6 -6 6 6
use M3_M2  M3_M2_96
timestamp 1543120812
transform 1 0 1448 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_97
timestamp 1543120812
transform 1 0 2808 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_98
timestamp 1543120812
transform 1 0 2776 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_99
timestamp 1543120812
transform 1 0 2504 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_100
timestamp 1543120812
transform 1 0 2360 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_101
timestamp 1543120812
transform 1 0 2984 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_102
timestamp 1543120812
transform 1 0 2968 0 1 2930
box -6 -6 6 6
use M3_M2  M3_M2_103
timestamp 1543120812
transform 1 0 2744 0 1 2090
box -6 -6 6 6
use M3_M2  M3_M2_104
timestamp 1543120812
transform 1 0 2744 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_105
timestamp 1543120812
transform 1 0 2632 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_106
timestamp 1543120812
transform 1 0 2632 0 1 2930
box -6 -6 6 6
use M3_M2  M3_M2_107
timestamp 1543120812
transform 1 0 2616 0 1 2090
box -6 -6 6 6
use M3_M2  M3_M2_108
timestamp 1543120812
transform 1 0 2568 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_109
timestamp 1543120812
transform 1 0 2520 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_110
timestamp 1543120812
transform 1 0 2392 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_111
timestamp 1543120812
transform 1 0 2360 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_112
timestamp 1543120812
transform 1 0 2312 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_113
timestamp 1543120812
transform 1 0 1960 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_114
timestamp 1543120812
transform 1 0 1832 0 1 3030
box -6 -6 6 6
use M3_M2  M3_M2_115
timestamp 1543120812
transform 1 0 1768 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_116
timestamp 1543120812
transform 1 0 1688 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_117
timestamp 1543120812
transform 1 0 1656 0 1 3030
box -6 -6 6 6
use M3_M2  M3_M2_118
timestamp 1543120812
transform 1 0 1656 0 1 2810
box -6 -6 6 6
use M3_M2  M3_M2_119
timestamp 1543120812
transform 1 0 1592 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_120
timestamp 1543120812
transform 1 0 1592 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_121
timestamp 1543120812
transform 1 0 1576 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_122
timestamp 1543120812
transform 1 0 1432 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_123
timestamp 1543120812
transform 1 0 1432 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_124
timestamp 1543120812
transform 1 0 1368 0 1 2810
box -6 -6 6 6
use M3_M2  M3_M2_125
timestamp 1543120812
transform 1 0 1352 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_126
timestamp 1543120812
transform 1 0 1336 0 1 3030
box -6 -6 6 6
use M3_M2  M3_M2_127
timestamp 1543120812
transform 1 0 1944 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_128
timestamp 1543120812
transform 1 0 1880 0 1 2550
box -6 -6 6 6
use M3_M2  M3_M2_129
timestamp 1543120812
transform 1 0 1880 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_130
timestamp 1543120812
transform 1 0 1784 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_131
timestamp 1543120812
transform 1 0 1720 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_132
timestamp 1543120812
transform 1 0 1672 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_133
timestamp 1543120812
transform 1 0 1640 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_134
timestamp 1543120812
transform 1 0 1640 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_135
timestamp 1543120812
transform 1 0 1608 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_136
timestamp 1543120812
transform 1 0 1608 0 1 2550
box -6 -6 6 6
use M3_M2  M3_M2_137
timestamp 1543120812
transform 1 0 1224 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_138
timestamp 1543120812
transform 1 0 2520 0 1 1070
box -6 -6 6 6
use M3_M2  M3_M2_139
timestamp 1543120812
transform 1 0 2472 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_140
timestamp 1543120812
transform 1 0 2472 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_141
timestamp 1543120812
transform 1 0 2408 0 1 2650
box -6 -6 6 6
use M3_M2  M3_M2_142
timestamp 1543120812
transform 1 0 2408 0 1 1070
box -6 -6 6 6
use M3_M2  M3_M2_143
timestamp 1543120812
transform 1 0 2280 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_144
timestamp 1543120812
transform 1 0 2264 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_145
timestamp 1543120812
transform 1 0 2216 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_146
timestamp 1543120812
transform 1 0 2200 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_147
timestamp 1543120812
transform 1 0 2200 0 1 1070
box -6 -6 6 6
use M3_M2  M3_M2_148
timestamp 1543120812
transform 1 0 2648 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_149
timestamp 1543120812
transform 1 0 2632 0 1 2650
box -6 -6 6 6
use M3_M2  M3_M2_150
timestamp 1543120812
transform 1 0 2472 0 1 2650
box -6 -6 6 6
use M3_M2  M3_M2_151
timestamp 1543120812
transform 1 0 2424 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_152
timestamp 1543120812
transform 1 0 2408 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_153
timestamp 1543120812
transform 1 0 2296 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_154
timestamp 1543120812
transform 1 0 2232 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_155
timestamp 1543120812
transform 1 0 1560 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_156
timestamp 1543120812
transform 1 0 1496 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_157
timestamp 1543120812
transform 1 0 1464 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_158
timestamp 1543120812
transform 1 0 1432 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_159
timestamp 1543120812
transform 1 0 1304 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_160
timestamp 1543120812
transform 1 0 1304 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_161
timestamp 1543120812
transform 1 0 1208 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_162
timestamp 1543120812
transform 1 0 1208 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_163
timestamp 1543120812
transform 1 0 1464 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_164
timestamp 1543120812
transform 1 0 1368 0 1 1730
box -6 -6 6 6
use M3_M2  M3_M2_165
timestamp 1543120812
transform 1 0 1336 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_166
timestamp 1543120812
transform 1 0 1224 0 1 2170
box -6 -6 6 6
use M3_M2  M3_M2_167
timestamp 1543120812
transform 1 0 1224 0 1 1730
box -6 -6 6 6
use M3_M2  M3_M2_168
timestamp 1543120812
transform 1 0 1016 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_169
timestamp 1543120812
transform 1 0 984 0 1 2170
box -6 -6 6 6
use M3_M2  M3_M2_170
timestamp 1543120812
transform 1 0 952 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_171
timestamp 1543120812
transform 1 0 2520 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_172
timestamp 1543120812
transform 1 0 2488 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_173
timestamp 1543120812
transform 1 0 2248 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_174
timestamp 1543120812
transform 1 0 2248 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_175
timestamp 1543120812
transform 1 0 2152 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_176
timestamp 1543120812
transform 1 0 2088 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_177
timestamp 1543120812
transform 1 0 2088 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_178
timestamp 1543120812
transform 1 0 2024 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_179
timestamp 1543120812
transform 1 0 2024 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_180
timestamp 1543120812
transform 1 0 2696 0 1 2650
box -6 -6 6 6
use M3_M2  M3_M2_181
timestamp 1543120812
transform 1 0 2632 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_182
timestamp 1543120812
transform 1 0 2632 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_183
timestamp 1543120812
transform 1 0 2360 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_184
timestamp 1543120812
transform 1 0 2328 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_185
timestamp 1543120812
transform 1 0 2232 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_186
timestamp 1543120812
transform 1 0 2200 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_187
timestamp 1543120812
transform 1 0 1640 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_188
timestamp 1543120812
transform 1 0 1544 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_189
timestamp 1543120812
transform 1 0 1528 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_190
timestamp 1543120812
transform 1 0 1512 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_191
timestamp 1543120812
transform 1 0 1176 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_192
timestamp 1543120812
transform 1 0 1176 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_193
timestamp 1543120812
transform 1 0 1032 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_194
timestamp 1543120812
transform 1 0 1032 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_195
timestamp 1543120812
transform 1 0 1400 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_196
timestamp 1543120812
transform 1 0 1400 0 1 2130
box -6 -6 6 6
use M3_M2  M3_M2_197
timestamp 1543120812
transform 1 0 1320 0 1 2130
box -6 -6 6 6
use M3_M2  M3_M2_198
timestamp 1543120812
transform 1 0 1256 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_199
timestamp 1543120812
transform 1 0 1048 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_200
timestamp 1543120812
transform 1 0 904 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_201
timestamp 1543120812
transform 1 0 904 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_202
timestamp 1543120812
transform 1 0 2744 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_203
timestamp 1543120812
transform 1 0 2520 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_204
timestamp 1543120812
transform 1 0 2504 0 1 2350
box -6 -6 6 6
use M3_M2  M3_M2_205
timestamp 1543120812
transform 1 0 2200 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_206
timestamp 1543120812
transform 1 0 2136 0 1 2350
box -6 -6 6 6
use M3_M2  M3_M2_207
timestamp 1543120812
transform 1 0 2040 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_208
timestamp 1543120812
transform 1 0 2616 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_209
timestamp 1543120812
transform 1 0 2312 0 1 2970
box -6 -6 6 6
use M3_M2  M3_M2_210
timestamp 1543120812
transform 1 0 2264 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_211
timestamp 1543120812
transform 1 0 2088 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_212
timestamp 1543120812
transform 1 0 2088 0 1 2970
box -6 -6 6 6
use M3_M2  M3_M2_213
timestamp 1543120812
transform 1 0 3160 0 1 3330
box -6 -6 6 6
use M3_M2  M3_M2_214
timestamp 1543120812
transform 1 0 2904 0 1 3330
box -6 -6 6 6
use M3_M2  M3_M2_215
timestamp 1543120812
transform 1 0 1720 0 1 3330
box -6 -6 6 6
use M3_M2  M3_M2_216
timestamp 1543120812
transform 1 0 1624 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_217
timestamp 1543120812
transform 1 0 1400 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_218
timestamp 1543120812
transform 1 0 2936 0 1 3290
box -6 -6 6 6
use M3_M2  M3_M2_219
timestamp 1543120812
transform 1 0 2712 0 1 3290
box -6 -6 6 6
use M3_M2  M3_M2_220
timestamp 1543120812
transform 1 0 2200 0 1 3290
box -6 -6 6 6
use M3_M2  M3_M2_221
timestamp 1543120812
transform 1 0 2200 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_222
timestamp 1543120812
transform 1 0 1624 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_223
timestamp 1543120812
transform 1 0 1352 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_224
timestamp 1543120812
transform 1 0 1336 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_225
timestamp 1543120812
transform 1 0 2232 0 1 3170
box -6 -6 6 6
use M3_M2  M3_M2_226
timestamp 1543120812
transform 1 0 2104 0 1 3170
box -6 -6 6 6
use M3_M2  M3_M2_227
timestamp 1543120812
transform 1 0 2104 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_228
timestamp 1543120812
transform 1 0 1928 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_229
timestamp 1543120812
transform 1 0 2984 0 1 2970
box -6 -6 6 6
use M3_M2  M3_M2_230
timestamp 1543120812
transform 1 0 2824 0 1 2970
box -6 -6 6 6
use M3_M2  M3_M2_231
timestamp 1543120812
transform 1 0 1464 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_232
timestamp 1543120812
transform 1 0 1240 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_233
timestamp 1543120812
transform 1 0 1352 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_234
timestamp 1543120812
transform 1 0 1128 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_235
timestamp 1543120812
transform 1 0 1032 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_236
timestamp 1543120812
transform 1 0 3144 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_237
timestamp 1543120812
transform 1 0 2920 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_238
timestamp 1543120812
transform 1 0 2712 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_239
timestamp 1543120812
transform 1 0 1224 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_240
timestamp 1543120812
transform 1 0 1112 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_241
timestamp 1543120812
transform 1 0 1144 0 1 2350
box -6 -6 6 6
use M3_M2  M3_M2_242
timestamp 1543120812
transform 1 0 968 0 1 2350
box -6 -6 6 6
use M3_M2  M3_M2_243
timestamp 1543120812
transform 1 0 1000 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_244
timestamp 1543120812
transform 1 0 872 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_245
timestamp 1543120812
transform 1 0 2760 0 1 590
box -6 -6 6 6
use M3_M2  M3_M2_246
timestamp 1543120812
transform 1 0 2616 0 1 590
box -6 -6 6 6
use M3_M2  M3_M2_247
timestamp 1543120812
transform 1 0 3672 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_248
timestamp 1543120812
transform 1 0 3368 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_249
timestamp 1543120812
transform 1 0 3400 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_250
timestamp 1543120812
transform 1 0 3240 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_251
timestamp 1543120812
transform 1 0 3448 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_252
timestamp 1543120812
transform 1 0 3384 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_253
timestamp 1543120812
transform 1 0 3560 0 1 1050
box -6 -6 6 6
use M3_M2  M3_M2_254
timestamp 1543120812
transform 1 0 3544 0 1 1170
box -6 -6 6 6
use M3_M2  M3_M2_255
timestamp 1543120812
transform 1 0 3576 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_256
timestamp 1543120812
transform 1 0 3528 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_257
timestamp 1543120812
transform 1 0 3352 0 1 670
box -6 -6 6 6
use M3_M2  M3_M2_258
timestamp 1543120812
transform 1 0 3304 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_259
timestamp 1543120812
transform 1 0 3496 0 1 430
box -6 -6 6 6
use M3_M2  M3_M2_260
timestamp 1543120812
transform 1 0 3096 0 1 430
box -6 -6 6 6
use M3_M2  M3_M2_261
timestamp 1543120812
transform 1 0 3320 0 1 370
box -6 -6 6 6
use M3_M2  M3_M2_262
timestamp 1543120812
transform 1 0 3224 0 1 370
box -6 -6 6 6
use M3_M2  M3_M2_263
timestamp 1543120812
transform 1 0 3224 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_264
timestamp 1543120812
transform 1 0 2952 0 1 370
box -6 -6 6 6
use M3_M2  M3_M2_265
timestamp 1543120812
transform 1 0 2920 0 1 350
box -6 -6 6 6
use M3_M2  M3_M2_266
timestamp 1543120812
transform 1 0 2536 0 1 350
box -6 -6 6 6
use M3_M2  M3_M2_267
timestamp 1543120812
transform 1 0 2840 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_268
timestamp 1543120812
transform 1 0 2424 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_269
timestamp 1543120812
transform 1 0 2616 0 1 610
box -6 -6 6 6
use M3_M2  M3_M2_270
timestamp 1543120812
transform 1 0 2504 0 1 610
box -6 -6 6 6
use M3_M2  M3_M2_271
timestamp 1543120812
transform 1 0 2344 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_272
timestamp 1543120812
transform 1 0 2184 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_273
timestamp 1543120812
transform 1 0 2392 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_274
timestamp 1543120812
transform 1 0 2232 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_275
timestamp 1543120812
transform 1 0 3560 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_276
timestamp 1543120812
transform 1 0 3496 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_277
timestamp 1543120812
transform 1 0 3448 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_278
timestamp 1543120812
transform 1 0 3384 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_279
timestamp 1543120812
transform 1 0 3288 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_280
timestamp 1543120812
transform 1 0 3592 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_281
timestamp 1543120812
transform 1 0 3336 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_282
timestamp 1543120812
transform 1 0 3624 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_283
timestamp 1543120812
transform 1 0 3448 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_284
timestamp 1543120812
transform 1 0 3512 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_285
timestamp 1543120812
transform 1 0 3336 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_286
timestamp 1543120812
transform 1 0 3272 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_287
timestamp 1543120812
transform 1 0 3016 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_288
timestamp 1543120812
transform 1 0 2904 0 1 390
box -6 -6 6 6
use M3_M2  M3_M2_289
timestamp 1543120812
transform 1 0 3080 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_290
timestamp 1543120812
transform 1 0 2984 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_291
timestamp 1543120812
transform 1 0 2824 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_292
timestamp 1543120812
transform 1 0 2648 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_293
timestamp 1543120812
transform 1 0 3064 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_294
timestamp 1543120812
transform 1 0 2968 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_295
timestamp 1543120812
transform 1 0 2872 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_296
timestamp 1543120812
transform 1 0 2728 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_297
timestamp 1543120812
transform 1 0 2632 0 1 570
box -6 -6 6 6
use M3_M2  M3_M2_298
timestamp 1543120812
transform 1 0 2568 0 1 570
box -6 -6 6 6
use M3_M2  M3_M2_299
timestamp 1543120812
transform 1 0 2536 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_300
timestamp 1543120812
transform 1 0 2344 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_301
timestamp 1543120812
transform 1 0 2168 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_302
timestamp 1543120812
transform 1 0 1896 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_303
timestamp 1543120812
transform 1 0 2664 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_304
timestamp 1543120812
transform 1 0 2584 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_305
timestamp 1543120812
transform 1 0 2296 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_306
timestamp 1543120812
transform 1 0 2120 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_307
timestamp 1543120812
transform 1 0 1224 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_308
timestamp 1543120812
transform 1 0 1192 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_309
timestamp 1543120812
transform 1 0 1128 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_310
timestamp 1543120812
transform 1 0 1128 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_311
timestamp 1543120812
transform 1 0 952 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_312
timestamp 1543120812
transform 1 0 664 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_313
timestamp 1543120812
transform 1 0 760 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_314
timestamp 1543120812
transform 1 0 632 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_315
timestamp 1543120812
transform 1 0 1048 0 1 1390
box -6 -6 6 6
use M3_M2  M3_M2_316
timestamp 1543120812
transform 1 0 488 0 1 1390
box -6 -6 6 6
use M3_M2  M3_M2_317
timestamp 1543120812
transform 1 0 2776 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_318
timestamp 1543120812
transform 1 0 2696 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_319
timestamp 1543120812
transform 1 0 2472 0 1 1550
box -6 -6 6 6
use M3_M2  M3_M2_320
timestamp 1543120812
transform 1 0 1784 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_321
timestamp 1543120812
transform 1 0 1704 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_322
timestamp 1543120812
transform 1 0 808 0 1 1430
box -6 -6 6 6
use M3_M2  M3_M2_323
timestamp 1543120812
transform 1 0 744 0 1 1430
box -6 -6 6 6
use M3_M2  M3_M2_324
timestamp 1543120812
transform 1 0 2104 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_325
timestamp 1543120812
transform 1 0 2024 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_326
timestamp 1543120812
transform 1 0 2136 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_327
timestamp 1543120812
transform 1 0 2008 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_328
timestamp 1543120812
transform 1 0 1336 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_329
timestamp 1543120812
transform 1 0 1288 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_330
timestamp 1543120812
transform 1 0 2360 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_331
timestamp 1543120812
transform 1 0 2088 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_332
timestamp 1543120812
transform 1 0 3128 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_333
timestamp 1543120812
transform 1 0 2968 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_334
timestamp 1543120812
transform 1 0 2648 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_335
timestamp 1543120812
transform 1 0 2120 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_336
timestamp 1543120812
transform 1 0 2104 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_337
timestamp 1543120812
transform 1 0 1992 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_338
timestamp 1543120812
transform 1 0 1624 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_339
timestamp 1543120812
transform 1 0 1496 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_340
timestamp 1543120812
transform 1 0 1240 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_341
timestamp 1543120812
transform 1 0 1240 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_342
timestamp 1543120812
transform 1 0 888 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_343
timestamp 1543120812
transform 1 0 616 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_344
timestamp 1543120812
transform 1 0 1560 0 1 2450
box -6 -6 6 6
use M3_M2  M3_M2_345
timestamp 1543120812
transform 1 0 1320 0 1 2450
box -6 -6 6 6
use M3_M2  M3_M2_346
timestamp 1543120812
transform 1 0 1160 0 1 2450
box -6 -6 6 6
use M3_M2  M3_M2_347
timestamp 1543120812
transform 1 0 984 0 1 2450
box -6 -6 6 6
use M3_M2  M3_M2_348
timestamp 1543120812
transform 1 0 712 0 1 2430
box -6 -6 6 6
use M3_M2  M3_M2_349
timestamp 1543120812
transform 1 0 3352 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_350
timestamp 1543120812
transform 1 0 3224 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_351
timestamp 1543120812
transform 1 0 2792 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_352
timestamp 1543120812
transform 1 0 2376 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_353
timestamp 1543120812
transform 1 0 2248 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_354
timestamp 1543120812
transform 1 0 2248 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_355
timestamp 1543120812
transform 1 0 2136 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_356
timestamp 1543120812
transform 1 0 2632 0 1 3390
box -6 -6 6 6
use M3_M2  M3_M2_357
timestamp 1543120812
transform 1 0 2504 0 1 3390
box -6 -6 6 6
use M3_M2  M3_M2_358
timestamp 1543120812
transform 1 0 680 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_359
timestamp 1543120812
transform 1 0 552 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_360
timestamp 1543120812
transform 1 0 3160 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_361
timestamp 1543120812
transform 1 0 2952 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_362
timestamp 1543120812
transform 1 0 2952 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_363
timestamp 1543120812
transform 1 0 2648 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_364
timestamp 1543120812
transform 1 0 2424 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_365
timestamp 1543120812
transform 1 0 968 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_366
timestamp 1543120812
transform 1 0 776 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_367
timestamp 1543120812
transform 1 0 1256 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_368
timestamp 1543120812
transform 1 0 1048 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_369
timestamp 1543120812
transform 1 0 3016 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_370
timestamp 1543120812
transform 1 0 2536 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_371
timestamp 1543120812
transform 1 0 2872 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_372
timestamp 1543120812
transform 1 0 2632 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_373
timestamp 1543120812
transform 1 0 2376 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_374
timestamp 1543120812
transform 1 0 1912 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_375
timestamp 1543120812
transform 1 0 1912 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_376
timestamp 1543120812
transform 1 0 1784 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_377
timestamp 1543120812
transform 1 0 1752 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_378
timestamp 1543120812
transform 1 0 1256 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_379
timestamp 1543120812
transform 1 0 1256 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_380
timestamp 1543120812
transform 1 0 824 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_381
timestamp 1543120812
transform 1 0 808 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_382
timestamp 1543120812
transform 1 0 712 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_383
timestamp 1543120812
transform 1 0 1672 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_384
timestamp 1543120812
transform 1 0 1432 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_385
timestamp 1543120812
transform 1 0 1208 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_386
timestamp 1543120812
transform 1 0 904 0 1 2030
box -6 -6 6 6
use M3_M2  M3_M2_387
timestamp 1543120812
transform 1 0 3272 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_388
timestamp 1543120812
transform 1 0 2968 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_389
timestamp 1543120812
transform 1 0 2760 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_390
timestamp 1543120812
transform 1 0 2552 0 1 2370
box -6 -6 6 6
use M3_M2  M3_M2_391
timestamp 1543120812
transform 1 0 1752 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_392
timestamp 1543120812
transform 1 0 1608 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_393
timestamp 1543120812
transform 1 0 2872 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_394
timestamp 1543120812
transform 1 0 2824 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_395
timestamp 1543120812
transform 1 0 2600 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_396
timestamp 1543120812
transform 1 0 2600 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_397
timestamp 1543120812
transform 1 0 2440 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_398
timestamp 1543120812
transform 1 0 2440 0 1 670
box -6 -6 6 6
use M3_M2  M3_M2_399
timestamp 1543120812
transform 1 0 2072 0 1 670
box -6 -6 6 6
use M3_M2  M3_M2_400
timestamp 1543120812
transform 1 0 1816 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_401
timestamp 1543120812
transform 1 0 1448 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_402
timestamp 1543120812
transform 1 0 1416 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_403
timestamp 1543120812
transform 1 0 1304 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_404
timestamp 1543120812
transform 1 0 1240 0 1 1350
box -6 -6 6 6
use M3_M2  M3_M2_405
timestamp 1543120812
transform 1 0 1112 0 1 1350
box -6 -6 6 6
use M3_M2  M3_M2_406
timestamp 1543120812
transform 1 0 872 0 1 1350
box -6 -6 6 6
use M3_M2  M3_M2_407
timestamp 1543120812
transform 1 0 2488 0 1 1730
box -6 -6 6 6
use M3_M2  M3_M2_408
timestamp 1543120812
transform 1 0 2360 0 1 1730
box -6 -6 6 6
use M3_M2  M3_M2_409
timestamp 1543120812
transform 1 0 1784 0 1 1730
box -6 -6 6 6
use M3_M2  M3_M2_410
timestamp 1543120812
transform 1 0 2280 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_411
timestamp 1543120812
transform 1 0 1896 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_412
timestamp 1543120812
transform 1 0 1768 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_413
timestamp 1543120812
transform 1 0 2264 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_414
timestamp 1543120812
transform 1 0 2088 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_415
timestamp 1543120812
transform 1 0 1960 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_416
timestamp 1543120812
transform 1 0 1544 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_417
timestamp 1543120812
transform 1 0 1272 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_418
timestamp 1543120812
transform 1 0 2136 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_419
timestamp 1543120812
transform 1 0 2056 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_420
timestamp 1543120812
transform 1 0 1800 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_421
timestamp 1543120812
transform 1 0 1624 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_422
timestamp 1543120812
transform 1 0 1432 0 1 1930
box -6 -6 6 6
use M3_M2  M3_M2_423
timestamp 1543120812
transform 1 0 2104 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_424
timestamp 1543120812
transform 1 0 1608 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_425
timestamp 1543120812
transform 1 0 1144 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_426
timestamp 1543120812
transform 1 0 1048 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_427
timestamp 1543120812
transform 1 0 904 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_428
timestamp 1543120812
transform 1 0 728 0 1 770
box -6 -6 6 6
use M3_M2  M3_M2_429
timestamp 1543120812
transform 1 0 1176 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_430
timestamp 1543120812
transform 1 0 792 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_431
timestamp 1543120812
transform 1 0 776 0 1 930
box -6 -6 6 6
use M3_M2  M3_M2_432
timestamp 1543120812
transform 1 0 456 0 1 930
box -6 -6 6 6
use M3_M2  M3_M2_433
timestamp 1543120812
transform 1 0 2040 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_434
timestamp 1543120812
transform 1 0 1960 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_435
timestamp 1543120812
transform 1 0 648 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_436
timestamp 1543120812
transform 1 0 584 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_437
timestamp 1543120812
transform 1 0 808 0 1 3030
box -6 -6 6 6
use M3_M2  M3_M2_438
timestamp 1543120812
transform 1 0 728 0 1 3030
box -6 -6 6 6
use M3_M2  M3_M2_439
timestamp 1543120812
transform 1 0 2536 0 1 3430
box -6 -6 6 6
use M3_M2  M3_M2_440
timestamp 1543120812
transform 1 0 2488 0 1 3430
box -6 -6 6 6
use M3_M2  M3_M2_441
timestamp 1543120812
transform 1 0 1752 0 1 270
box -6 -6 6 6
use M3_M2  M3_M2_442
timestamp 1543120812
transform 1 0 1480 0 1 270
box -6 -6 6 6
use M3_M2  M3_M2_443
timestamp 1543120812
transform 1 0 2616 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_444
timestamp 1543120812
transform 1 0 2360 0 1 1150
box -6 -6 6 6
use M3_M2  M3_M2_445
timestamp 1543120812
transform 1 0 2280 0 1 1870
box -6 -6 6 6
use M3_M2  M3_M2_446
timestamp 1543120812
transform 1 0 2200 0 1 1150
box -6 -6 6 6
use M3_M2  M3_M2_447
timestamp 1543120812
transform 1 0 1816 0 1 1870
box -6 -6 6 6
use M3_M2  M3_M2_448
timestamp 1543120812
transform 1 0 1816 0 1 1670
box -6 -6 6 6
use M3_M2  M3_M2_449
timestamp 1543120812
transform 1 0 1800 0 1 1150
box -6 -6 6 6
use M3_M2  M3_M2_450
timestamp 1543120812
transform 1 0 1720 0 1 450
box -6 -6 6 6
use M3_M2  M3_M2_451
timestamp 1543120812
transform 1 0 1688 0 1 1150
box -6 -6 6 6
use M3_M2  M3_M2_452
timestamp 1543120812
transform 1 0 1464 0 1 1670
box -6 -6 6 6
use M3_M2  M3_M2_453
timestamp 1543120812
transform 1 0 1304 0 1 1670
box -6 -6 6 6
use M3_M2  M3_M2_454
timestamp 1543120812
transform 1 0 1176 0 1 430
box -6 -6 6 6
use M3_M2  M3_M2_455
timestamp 1543120812
transform 1 0 680 0 1 590
box -6 -6 6 6
use M3_M2  M3_M2_456
timestamp 1543120812
transform 1 0 680 0 1 430
box -6 -6 6 6
use M3_M2  M3_M2_457
timestamp 1543120812
transform 1 0 344 0 1 590
box -6 -6 6 6
use M3_M2  M3_M2_458
timestamp 1543120812
transform 1 0 3064 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_459
timestamp 1543120812
transform 1 0 3000 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_460
timestamp 1543120812
transform 1 0 2968 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_461
timestamp 1543120812
transform 1 0 2856 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_462
timestamp 1543120812
transform 1 0 2776 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_463
timestamp 1543120812
transform 1 0 2776 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_464
timestamp 1543120812
transform 1 0 2728 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_465
timestamp 1543120812
transform 1 0 2552 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_466
timestamp 1543120812
transform 1 0 2552 0 1 750
box -6 -6 6 6
use M3_M2  M3_M2_467
timestamp 1543120812
transform 1 0 2360 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_468
timestamp 1543120812
transform 1 0 2184 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_469
timestamp 1543120812
transform 1 0 1896 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_470
timestamp 1543120812
transform 1 0 1864 0 1 370
box -6 -6 6 6
use M3_M2  M3_M2_471
timestamp 1543120812
transform 1 0 1672 0 1 370
box -6 -6 6 6
use M3_M2  M3_M2_472
timestamp 1543120812
transform 1 0 3320 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_473
timestamp 1543120812
transform 1 0 3272 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_474
timestamp 1543120812
transform 1 0 3240 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_475
timestamp 1543120812
transform 1 0 3144 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_476
timestamp 1543120812
transform 1 0 3096 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_477
timestamp 1543120812
transform 1 0 3000 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_478
timestamp 1543120812
transform 1 0 2856 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_479
timestamp 1543120812
transform 1 0 2840 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_480
timestamp 1543120812
transform 1 0 2536 0 1 3470
box -6 -6 6 6
use M3_M2  M3_M2_481
timestamp 1543120812
transform 1 0 2168 0 1 3470
box -6 -6 6 6
use M3_M2  M3_M2_482
timestamp 1543120812
transform 1 0 1208 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_483
timestamp 1543120812
transform 1 0 936 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_484
timestamp 1543120812
transform 1 0 824 0 1 3490
box -6 -6 6 6
use M3_M2  M3_M2_485
timestamp 1543120812
transform 1 0 744 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_486
timestamp 1543120812
transform 1 0 3176 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_487
timestamp 1543120812
transform 1 0 3160 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_488
timestamp 1543120812
transform 1 0 3080 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_489
timestamp 1543120812
transform 1 0 3032 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_490
timestamp 1543120812
transform 1 0 2744 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_491
timestamp 1543120812
transform 1 0 2488 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_492
timestamp 1543120812
transform 1 0 1976 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_493
timestamp 1543120812
transform 1 0 1144 0 1 3450
box -6 -6 6 6
use M3_M2  M3_M2_494
timestamp 1543120812
transform 1 0 856 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_495
timestamp 1543120812
transform 1 0 760 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_496
timestamp 1543120812
transform 1 0 696 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_497
timestamp 1543120812
transform 1 0 600 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_498
timestamp 1543120812
transform 1 0 584 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_499
timestamp 1543120812
transform 1 0 3160 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_500
timestamp 1543120812
transform 1 0 3160 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_501
timestamp 1543120812
transform 1 0 3080 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_502
timestamp 1543120812
transform 1 0 3000 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_503
timestamp 1543120812
transform 1 0 2968 0 1 2950
box -6 -6 6 6
use M3_M2  M3_M2_504
timestamp 1543120812
transform 1 0 2936 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_505
timestamp 1543120812
transform 1 0 2824 0 1 2950
box -6 -6 6 6
use M3_M2  M3_M2_506
timestamp 1543120812
transform 1 0 2824 0 1 2710
box -6 -6 6 6
use M3_M2  M3_M2_507
timestamp 1543120812
transform 1 0 2776 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_508
timestamp 1543120812
transform 1 0 2680 0 1 2190
box -6 -6 6 6
use M3_M2  M3_M2_509
timestamp 1543120812
transform 1 0 2440 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_510
timestamp 1543120812
transform 1 0 2056 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_511
timestamp 1543120812
transform 1 0 1640 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_512
timestamp 1543120812
transform 1 0 1448 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_513
timestamp 1543120812
transform 1 0 1384 0 1 1330
box -6 -6 6 6
use M3_M2  M3_M2_514
timestamp 1543120812
transform 1 0 1384 0 1 710
box -6 -6 6 6
use M3_M2  M3_M2_515
timestamp 1543120812
transform 1 0 1080 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_516
timestamp 1543120812
transform 1 0 1080 0 1 1330
box -6 -6 6 6
use M3_M2  M3_M2_517
timestamp 1543120812
transform 1 0 968 0 1 2150
box -6 -6 6 6
use M3_M2  M3_M2_518
timestamp 1543120812
transform 1 0 840 0 1 3170
box -6 -6 6 6
use M3_M2  M3_M2_519
timestamp 1543120812
transform 1 0 840 0 1 2150
box -6 -6 6 6
use M3_M2  M3_M2_520
timestamp 1543120812
transform 1 0 808 0 1 2570
box -6 -6 6 6
use M3_M2  M3_M2_521
timestamp 1543120812
transform 1 0 808 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_522
timestamp 1543120812
transform 1 0 696 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_523
timestamp 1543120812
transform 1 0 616 0 1 2310
box -6 -6 6 6
use M3_M2  M3_M2_524
timestamp 1543120812
transform 1 0 3480 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_525
timestamp 1543120812
transform 1 0 3368 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_526
timestamp 1543120812
transform 1 0 3480 0 1 1810
box -6 -6 6 6
use M3_M2  M3_M2_527
timestamp 1543120812
transform 1 0 3368 0 1 1810
box -6 -6 6 6
use M3_M2  M3_M2_528
timestamp 1543120812
transform 1 0 2952 0 1 810
box -6 -6 6 6
use M3_M2  M3_M2_529
timestamp 1543120812
transform 1 0 2824 0 1 810
box -6 -6 6 6
use M3_M2  M3_M2_530
timestamp 1543120812
transform 1 0 3208 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_531
timestamp 1543120812
transform 1 0 3080 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_532
timestamp 1543120812
transform 1 0 3192 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_533
timestamp 1543120812
transform 1 0 3064 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_534
timestamp 1543120812
transform 1 0 3080 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_535
timestamp 1543120812
transform 1 0 2952 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_536
timestamp 1543120812
transform 1 0 2024 0 1 410
box -6 -6 6 6
use M3_M2  M3_M2_537
timestamp 1543120812
transform 1 0 1928 0 1 410
box -6 -6 6 6
use M3_M2  M3_M2_538
timestamp 1543120812
transform 1 0 2728 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_539
timestamp 1543120812
transform 1 0 2616 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_540
timestamp 1543120812
transform 1 0 3048 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_541
timestamp 1543120812
transform 1 0 2888 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_542
timestamp 1543120812
transform 1 0 1912 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_543
timestamp 1543120812
transform 1 0 1736 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_544
timestamp 1543120812
transform 1 0 1912 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_545
timestamp 1543120812
transform 1 0 1848 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_546
timestamp 1543120812
transform 1 0 2024 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_547
timestamp 1543120812
transform 1 0 2008 0 1 3310
box -6 -6 6 6
use M3_M2  M3_M2_548
timestamp 1543120812
transform 1 0 1864 0 1 3310
box -6 -6 6 6
use M3_M2  M3_M2_549
timestamp 1543120812
transform 1 0 1864 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_550
timestamp 1543120812
transform 1 0 1944 0 1 3410
box -6 -6 6 6
use M3_M2  M3_M2_551
timestamp 1543120812
transform 1 0 1800 0 1 3410
box -6 -6 6 6
use M3_M2  M3_M2_552
timestamp 1543120812
transform 1 0 1608 0 1 3410
box -6 -6 6 6
use M3_M2  M3_M2_553
timestamp 1543120812
transform 1 0 792 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_554
timestamp 1543120812
transform 1 0 568 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_555
timestamp 1543120812
transform 1 0 424 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_556
timestamp 1543120812
transform 1 0 616 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_557
timestamp 1543120812
transform 1 0 616 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_558
timestamp 1543120812
transform 1 0 408 0 1 3250
box -6 -6 6 6
use M3_M2  M3_M2_559
timestamp 1543120812
transform 1 0 408 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_560
timestamp 1543120812
transform 1 0 2072 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_561
timestamp 1543120812
transform 1 0 1928 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_562
timestamp 1543120812
transform 1 0 1560 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_563
timestamp 1543120812
transform 1 0 1240 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_564
timestamp 1543120812
transform 1 0 1240 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_565
timestamp 1543120812
transform 1 0 1128 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_566
timestamp 1543120812
transform 1 0 1768 0 1 1810
box -6 -6 6 6
use M3_M2  M3_M2_567
timestamp 1543120812
transform 1 0 1752 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_568
timestamp 1543120812
transform 1 0 1608 0 1 1810
box -6 -6 6 6
use M3_M2  M3_M2_569
timestamp 1543120812
transform 1 0 1592 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_570
timestamp 1543120812
transform 1 0 1592 0 1 1250
box -6 -6 6 6
use M3_M2  M3_M2_571
timestamp 1543120812
transform 1 0 1528 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_572
timestamp 1543120812
transform 1 0 1768 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_573
timestamp 1543120812
transform 1 0 1752 0 1 950
box -6 -6 6 6
use M3_M2  M3_M2_574
timestamp 1543120812
transform 1 0 1640 0 1 950
box -6 -6 6 6
use M3_M2  M3_M2_575
timestamp 1543120812
transform 1 0 1608 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_576
timestamp 1543120812
transform 1 0 1336 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_577
timestamp 1543120812
transform 1 0 1240 0 1 1690
box -6 -6 6 6
use M3_M2  M3_M2_578
timestamp 1543120812
transform 1 0 2472 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_579
timestamp 1543120812
transform 1 0 2328 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_580
timestamp 1543120812
transform 1 0 2264 0 1 930
box -6 -6 6 6
use M3_M2  M3_M2_581
timestamp 1543120812
transform 1 0 2152 0 1 930
box -6 -6 6 6
use M3_M2  M3_M2_582
timestamp 1543120812
transform 1 0 2072 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_583
timestamp 1543120812
transform 1 0 2184 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_584
timestamp 1543120812
transform 1 0 2040 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_585
timestamp 1543120812
transform 1 0 1992 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_586
timestamp 1543120812
transform 1 0 1496 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_587
timestamp 1543120812
transform 1 0 1304 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_588
timestamp 1543120812
transform 1 0 1208 0 1 1610
box -6 -6 6 6
use M3_M2  M3_M2_589
timestamp 1543120812
transform 1 0 2504 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_590
timestamp 1543120812
transform 1 0 2344 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_591
timestamp 1543120812
transform 1 0 2344 0 1 1330
box -6 -6 6 6
use M3_M2  M3_M2_592
timestamp 1543120812
transform 1 0 2264 0 1 1330
box -6 -6 6 6
use M3_M2  M3_M2_593
timestamp 1543120812
transform 1 0 2248 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_594
timestamp 1543120812
transform 1 0 2120 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_595
timestamp 1543120812
transform 1 0 1480 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_596
timestamp 1543120812
transform 1 0 1336 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_597
timestamp 1543120812
transform 1 0 1256 0 1 1070
box -6 -6 6 6
use M3_M2  M3_M2_598
timestamp 1543120812
transform 1 0 1160 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_599
timestamp 1543120812
transform 1 0 2232 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_600
timestamp 1543120812
transform 1 0 1928 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_601
timestamp 1543120812
transform 1 0 1720 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_602
timestamp 1543120812
transform 1 0 2472 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_603
timestamp 1543120812
transform 1 0 2392 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_604
timestamp 1543120812
transform 1 0 1736 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_605
timestamp 1543120812
transform 1 0 1192 0 1 1650
box -6 -6 6 6
use M3_M2  M3_M2_606
timestamp 1543120812
transform 1 0 984 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_607
timestamp 1543120812
transform 1 0 856 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_608
timestamp 1543120812
transform 1 0 872 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_609
timestamp 1543120812
transform 1 0 760 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_610
timestamp 1543120812
transform 1 0 760 0 1 1190
box -6 -6 6 6
use M3_M2  M3_M2_611
timestamp 1543120812
transform 1 0 632 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_612
timestamp 1543120812
transform 1 0 568 0 1 1630
box -6 -6 6 6
use M3_M2  M3_M2_613
timestamp 1543120812
transform 1 0 904 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_614
timestamp 1543120812
transform 1 0 600 0 1 1530
box -6 -6 6 6
use M3_M2  M3_M2_615
timestamp 1543120812
transform 1 0 760 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_616
timestamp 1543120812
transform 1 0 600 0 1 850
box -6 -6 6 6
use M3_M2  M3_M2_617
timestamp 1543120812
transform 1 0 808 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_618
timestamp 1543120812
transform 1 0 472 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_619
timestamp 1543120812
transform 1 0 936 0 1 570
box -6 -6 6 6
use M3_M2  M3_M2_620
timestamp 1543120812
transform 1 0 728 0 1 570
box -6 -6 6 6
use M3_M2  M3_M2_621
timestamp 1543120812
transform 1 0 1016 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_622
timestamp 1543120812
transform 1 0 744 0 1 1090
box -6 -6 6 6
use M3_M2  M3_M2_623
timestamp 1543120812
transform 1 0 824 0 1 1050
box -6 -6 6 6
use M3_M2  M3_M2_624
timestamp 1543120812
transform 1 0 728 0 1 1050
box -6 -6 6 6
use M3_M2  M3_M2_625
timestamp 1543120812
transform 1 0 1368 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_626
timestamp 1543120812
transform 1 0 1176 0 1 790
box -6 -6 6 6
use M3_M2  M3_M2_627
timestamp 1543120812
transform 1 0 1160 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_628
timestamp 1543120812
transform 1 0 968 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_629
timestamp 1543120812
transform 1 0 840 0 1 1130
box -6 -6 6 6
use M3_M2  M3_M2_630
timestamp 1543120812
transform 1 0 1272 0 1 1470
box -6 -6 6 6
use M3_M2  M3_M2_631
timestamp 1543120812
transform 1 0 968 0 1 1470
box -6 -6 6 6
use M3_M2  M3_M2_632
timestamp 1543120812
transform 1 0 776 0 1 1470
box -6 -6 6 6
use M3_M2  M3_M2_633
timestamp 1543120812
transform 1 0 1192 0 1 830
box -6 -6 6 6
use M3_M2  M3_M2_634
timestamp 1543120812
transform 1 0 952 0 1 830
box -6 -6 6 6
use M3_M2  M3_M2_635
timestamp 1543120812
transform 1 0 1800 0 1 1370
box -6 -6 6 6
use M3_M2  M3_M2_636
timestamp 1543120812
transform 1 0 1160 0 1 1370
box -6 -6 6 6
use M3_M2  M3_M2_637
timestamp 1543120812
transform 1 0 1016 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_638
timestamp 1543120812
transform 1 0 968 0 1 1230
box -6 -6 6 6
use M3_M2  M3_M2_639
timestamp 1543120812
transform 1 0 1928 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_640
timestamp 1543120812
transform 1 0 1240 0 1 1490
box -6 -6 6 6
use M3_M2  M3_M2_641
timestamp 1543120812
transform 1 0 1416 0 1 1410
box -6 -6 6 6
use M3_M2  M3_M2_642
timestamp 1543120812
transform 1 0 1256 0 1 1410
box -6 -6 6 6
use M3_M2  M3_M2_643
timestamp 1543120812
transform 1 0 1960 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_644
timestamp 1543120812
transform 1 0 1480 0 1 990
box -6 -6 6 6
use M3_M2  M3_M2_645
timestamp 1543120812
transform 1 0 2088 0 1 1050
box -6 -6 6 6
use M3_M2  M3_M2_646
timestamp 1543120812
transform 1 0 1992 0 1 1050
box -6 -6 6 6
use M3_M2  M3_M2_647
timestamp 1543120812
transform 1 0 2568 0 1 1430
box -6 -6 6 6
use M3_M2  M3_M2_648
timestamp 1543120812
transform 1 0 1784 0 1 1430
box -6 -6 6 6
use M3_M2  M3_M2_649
timestamp 1543120812
transform 1 0 1528 0 1 1450
box -6 -6 6 6
use M3_M2  M3_M2_650
timestamp 1543120812
transform 1 0 1432 0 1 1450
box -6 -6 6 6
use M3_M2  M3_M2_651
timestamp 1543120812
transform 1 0 2200 0 1 1370
box -6 -6 6 6
use M3_M2  M3_M2_652
timestamp 1543120812
transform 1 0 1976 0 1 1370
box -6 -6 6 6
use M3_M2  M3_M2_653
timestamp 1543120812
transform 1 0 456 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_654
timestamp 1543120812
transform 1 0 392 0 1 3090
box -6 -6 6 6
use M3_M2  M3_M2_655
timestamp 1543120812
transform 1 0 1640 0 1 3570
box -6 -6 6 6
use M3_M2  M3_M2_656
timestamp 1543120812
transform 1 0 1480 0 1 3570
box -6 -6 6 6
use M3_M2  M3_M2_657
timestamp 1543120812
transform 1 0 1880 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_658
timestamp 1543120812
transform 1 0 1704 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_659
timestamp 1543120812
transform 1 0 2168 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_660
timestamp 1543120812
transform 1 0 1736 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_661
timestamp 1543120812
transform 1 0 2536 0 1 2570
box -6 -6 6 6
use M3_M2  M3_M2_662
timestamp 1543120812
transform 1 0 1752 0 1 2570
box -6 -6 6 6
use M3_M2  M3_M2_663
timestamp 1543120812
transform 1 0 1800 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_664
timestamp 1543120812
transform 1 0 1224 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_665
timestamp 1543120812
transform 1 0 2776 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_666
timestamp 1543120812
transform 1 0 1816 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_667
timestamp 1543120812
transform 1 0 2792 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_668
timestamp 1543120812
transform 1 0 2648 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_669
timestamp 1543120812
transform 1 0 1192 0 1 2810
box -6 -6 6 6
use M3_M2  M3_M2_670
timestamp 1543120812
transform 1 0 1032 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_671
timestamp 1543120812
transform 1 0 1544 0 1 2270
box -6 -6 6 6
use M3_M2  M3_M2_672
timestamp 1543120812
transform 1 0 1416 0 1 2270
box -6 -6 6 6
use M3_M2  M3_M2_673
timestamp 1543120812
transform 1 0 1672 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_674
timestamp 1543120812
transform 1 0 1368 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_675
timestamp 1543120812
transform 1 0 1816 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_676
timestamp 1543120812
transform 1 0 1528 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_677
timestamp 1543120812
transform 1 0 1912 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_678
timestamp 1543120812
transform 1 0 1864 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_679
timestamp 1543120812
transform 1 0 1816 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_680
timestamp 1543120812
transform 1 0 1368 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_681
timestamp 1543120812
transform 1 0 1928 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_682
timestamp 1543120812
transform 1 0 1224 0 1 2730
box -6 -6 6 6
use M3_M2  M3_M2_683
timestamp 1543120812
transform 1 0 2504 0 1 2690
box -6 -6 6 6
use M3_M2  M3_M2_684
timestamp 1543120812
transform 1 0 1864 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_685
timestamp 1543120812
transform 1 0 2488 0 1 2770
box -6 -6 6 6
use M3_M2  M3_M2_686
timestamp 1543120812
transform 1 0 2472 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_687
timestamp 1543120812
transform 1 0 1240 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_688
timestamp 1543120812
transform 1 0 920 0 1 2870
box -6 -6 6 6
use M3_M2  M3_M2_689
timestamp 1543120812
transform 1 0 2056 0 1 2530
box -6 -6 6 6
use M3_M2  M3_M2_690
timestamp 1543120812
transform 1 0 1944 0 1 2530
box -6 -6 6 6
use M3_M2  M3_M2_691
timestamp 1543120812
transform 1 0 2440 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_692
timestamp 1543120812
transform 1 0 1992 0 1 2630
box -6 -6 6 6
use M3_M2  M3_M2_693
timestamp 1543120812
transform 1 0 1448 0 1 2650
box -6 -6 6 6
use M3_M2  M3_M2_694
timestamp 1543120812
transform 1 0 1384 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_695
timestamp 1543120812
transform 1 0 2344 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_696
timestamp 1543120812
transform 1 0 1896 0 1 2810
box -6 -6 6 6
use M3_M2  M3_M2_697
timestamp 1543120812
transform 1 0 2232 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_698
timestamp 1543120812
transform 1 0 1992 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_699
timestamp 1543120812
transform 1 0 2024 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_700
timestamp 1543120812
transform 1 0 2008 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_701
timestamp 1543120812
transform 1 0 1832 0 1 2890
box -6 -6 6 6
use M3_M2  M3_M2_702
timestamp 1543120812
transform 1 0 1832 0 1 2830
box -6 -6 6 6
use M3_M2  M3_M2_703
timestamp 1543120812
transform 1 0 1832 0 1 2790
box -6 -6 6 6
use M3_M2  M3_M2_704
timestamp 1543120812
transform 1 0 1832 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_705
timestamp 1543120812
transform 1 0 1928 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_706
timestamp 1543120812
transform 1 0 1544 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_707
timestamp 1543120812
transform 1 0 2248 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_708
timestamp 1543120812
transform 1 0 1992 0 1 2330
box -6 -6 6 6
use M3_M2  M3_M2_709
timestamp 1543120812
transform 1 0 2040 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_710
timestamp 1543120812
transform 1 0 1960 0 1 2250
box -6 -6 6 6
use M3_M2  M3_M2_711
timestamp 1543120812
transform 1 0 2440 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_712
timestamp 1543120812
transform 1 0 2344 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_713
timestamp 1543120812
transform 1 0 2584 0 1 2170
box -6 -6 6 6
use M3_M2  M3_M2_714
timestamp 1543120812
transform 1 0 2360 0 1 2170
box -6 -6 6 6
use M3_M2  M3_M2_715
timestamp 1543120812
transform 1 0 1928 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_716
timestamp 1543120812
transform 1 0 1784 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_717
timestamp 1543120812
transform 1 0 1576 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_718
timestamp 1543120812
transform 1 0 1496 0 1 2590
box -6 -6 6 6
use M3_M2  M3_M2_719
timestamp 1543120812
transform 1 0 1880 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_720
timestamp 1543120812
transform 1 0 1736 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_721
timestamp 1543120812
transform 1 0 2648 0 1 3130
box -6 -6 6 6
use M3_M2  M3_M2_722
timestamp 1543120812
transform 1 0 1896 0 1 3130
box -6 -6 6 6
use M3_M2  M3_M2_723
timestamp 1543120812
transform 1 0 1912 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_724
timestamp 1543120812
transform 1 0 1592 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_725
timestamp 1543120812
transform 1 0 1944 0 1 2910
box -6 -6 6 6
use M3_M2  M3_M2_726
timestamp 1543120812
transform 1 0 1784 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_727
timestamp 1543120812
transform 1 0 1720 0 1 2910
box -6 -6 6 6
use M3_M2  M3_M2_728
timestamp 1543120812
transform 1 0 1720 0 1 2670
box -6 -6 6 6
use M3_M2  M3_M2_729
timestamp 1543120812
transform 1 0 2776 0 1 2510
box -6 -6 6 6
use M3_M2  M3_M2_730
timestamp 1543120812
transform 1 0 1848 0 1 2510
box -6 -6 6 6
use M3_M2  M3_M2_731
timestamp 1543120812
transform 1 0 2728 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_732
timestamp 1543120812
transform 1 0 1960 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_733
timestamp 1543120812
transform 1 0 1896 0 1 2230
box -6 -6 6 6
use M3_M2  M3_M2_734
timestamp 1543120812
transform 1 0 1752 0 1 2230
box -6 -6 6 6
use M3_M2  M3_M2_735
timestamp 1543120812
transform 1 0 1608 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_736
timestamp 1543120812
transform 1 0 1464 0 1 3010
box -6 -6 6 6
use M3_M2  M3_M2_737
timestamp 1543120812
transform 1 0 2872 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_738
timestamp 1543120812
transform 1 0 2664 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_739
timestamp 1543120812
transform 1 0 920 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_740
timestamp 1543120812
transform 1 0 712 0 1 3230
box -6 -6 6 6
use M3_M2  M3_M2_741
timestamp 1543120812
transform 1 0 1528 0 1 3270
box -6 -6 6 6
use M3_M2  M3_M2_742
timestamp 1543120812
transform 1 0 696 0 1 3270
box -6 -6 6 6
use M3_M2  M3_M2_743
timestamp 1543120812
transform 1 0 1048 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_744
timestamp 1543120812
transform 1 0 984 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_745
timestamp 1543120812
transform 1 0 872 0 1 2390
box -6 -6 6 6
use M3_M2  M3_M2_746
timestamp 1543120812
transform 1 0 856 0 1 3190
box -6 -6 6 6
use M3_M2  M3_M2_747
timestamp 1543120812
transform 1 0 1112 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_748
timestamp 1543120812
transform 1 0 1016 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_749
timestamp 1543120812
transform 1 0 808 0 1 3150
box -6 -6 6 6
use M3_M2  M3_M2_750
timestamp 1543120812
transform 1 0 1064 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_751
timestamp 1543120812
transform 1 0 552 0 1 2750
box -6 -6 6 6
use M3_M2  M3_M2_752
timestamp 1543120812
transform 1 0 1288 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_753
timestamp 1543120812
transform 1 0 1064 0 1 3050
box -6 -6 6 6
use M3_M2  M3_M2_754
timestamp 1543120812
transform 1 0 1192 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_755
timestamp 1543120812
transform 1 0 1064 0 1 2990
box -6 -6 6 6
use M3_M2  M3_M2_756
timestamp 1543120812
transform 1 0 2488 0 1 2930
box -6 -6 6 6
use M3_M2  M3_M2_757
timestamp 1543120812
transform 1 0 1096 0 1 2930
box -6 -6 6 6
use M3_M2  M3_M2_758
timestamp 1543120812
transform 1 0 1176 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_759
timestamp 1543120812
transform 1 0 1016 0 1 2210
box -6 -6 6 6
use M3_M2  M3_M2_760
timestamp 1543120812
transform 1 0 2520 0 1 2070
box -6 -6 6 6
use M3_M2  M3_M2_761
timestamp 1543120812
transform 1 0 1032 0 1 2070
box -6 -6 6 6
use M3_M2  M3_M2_762
timestamp 1543120812
transform 1 0 2392 0 1 3370
box -6 -6 6 6
use M3_M2  M3_M2_763
timestamp 1543120812
transform 1 0 1480 0 1 3370
box -6 -6 6 6
use M3_M2  M3_M2_764
timestamp 1543120812
transform 1 0 2712 0 1 3270
box -6 -6 6 6
use M3_M2  M3_M2_765
timestamp 1543120812
transform 1 0 2408 0 1 3270
box -6 -6 6 6
use M3_M2  M3_M2_766
timestamp 1543120812
transform 1 0 1096 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_767
timestamp 1543120812
transform 1 0 1016 0 1 2610
box -6 -6 6 6
use M3_M2  M3_M2_768
timestamp 1543120812
transform 1 0 2232 0 1 2490
box -6 -6 6 6
use M3_M2  M3_M2_769
timestamp 1543120812
transform 1 0 1064 0 1 2490
box -6 -6 6 6
use M3_M2  M3_M2_770
timestamp 1543120812
transform 1 0 3128 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_771
timestamp 1543120812
transform 1 0 2984 0 1 2290
box -6 -6 6 6
use M3_M2  M3_M2_772
timestamp 1543120812
transform 1 0 1016 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_773
timestamp 1543120812
transform 1 0 904 0 1 1970
box -6 -6 6 6
use M3_M2  M3_M2_774
timestamp 1543120812
transform 1 0 2968 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_775
timestamp 1543120812
transform 1 0 2776 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_776
timestamp 1543120812
transform 1 0 3064 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_777
timestamp 1543120812
transform 1 0 2920 0 1 2850
box -6 -6 6 6
use M3_M2  M3_M2_778
timestamp 1543120812
transform 1 0 904 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_779
timestamp 1543120812
transform 1 0 808 0 1 3070
box -6 -6 6 6
use M3_M2  M3_M2_780
timestamp 1543120812
transform 1 0 3192 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_781
timestamp 1543120812
transform 1 0 3080 0 1 3110
box -6 -6 6 6
use M3_M2  M3_M2_782
timestamp 1543120812
transform 1 0 856 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_783
timestamp 1543120812
transform 1 0 728 0 1 2410
box -6 -6 6 6
use M3_M2  M3_M2_784
timestamp 1543120812
transform 1 0 2216 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_785
timestamp 1543120812
transform 1 0 2104 0 1 2050
box -6 -6 6 6
use M3_M2  M3_M2_786
timestamp 1543120812
transform 1 0 1576 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_787
timestamp 1543120812
transform 1 0 1480 0 1 2010
box -6 -6 6 6
use M3_M2  M3_M2_788
timestamp 1543120812
transform 1 0 1224 0 1 1670
box -6 -6 6 6
use M3_M2  M3_M2_789
timestamp 1543120812
transform 1 0 1144 0 1 1670
box -6 -6 6 6
use M3_M2  M3_M2_790
timestamp 1543120812
transform 1 0 2424 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_791
timestamp 1543120812
transform 1 0 2248 0 1 1030
box -6 -6 6 6
use M3_M2  M3_M2_792
timestamp 1543120812
transform 1 0 1848 0 1 1270
box -6 -6 6 6
use M3_M2  M3_M2_793
timestamp 1543120812
transform 1 0 1736 0 1 1270
box -6 -6 6 6
use M3_M2  M3_M2_794
timestamp 1543120812
transform 1 0 1752 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_795
timestamp 1543120812
transform 1 0 1560 0 1 1830
box -6 -6 6 6
use M3_M2  M3_M2_796
timestamp 1543120812
transform 1 0 1864 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_797
timestamp 1543120812
transform 1 0 1752 0 1 1570
box -6 -6 6 6
use M3_M2  M3_M2_798
timestamp 1543120812
transform 1 0 2664 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_799
timestamp 1543120812
transform 1 0 2456 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_800
timestamp 1543120812
transform 1 0 2632 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_801
timestamp 1543120812
transform 1 0 2504 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_802
timestamp 1543120812
transform 1 0 568 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_803
timestamp 1543120812
transform 1 0 440 0 1 1110
box -6 -6 6 6
use M3_M2  M3_M2_804
timestamp 1543120812
transform 1 0 2424 0 1 1290
box -6 -6 6 6
use M3_M2  M3_M2_805
timestamp 1543120812
transform 1 0 2248 0 1 1290
box -6 -6 6 6
use M3_M2  M3_M2_806
timestamp 1543120812
transform 1 0 1512 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_807
timestamp 1543120812
transform 1 0 1336 0 1 290
box -6 -6 6 6
use M3_M2  M3_M2_808
timestamp 1543120812
transform 1 0 3176 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_809
timestamp 1543120812
transform 1 0 3112 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_810
timestamp 1543120812
transform 1 0 3112 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_811
timestamp 1543120812
transform 1 0 3016 0 1 1590
box -6 -6 6 6
use M3_M2  M3_M2_812
timestamp 1543120812
transform 1 0 2920 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_813
timestamp 1543120812
transform 1 0 2856 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_814
timestamp 1543120812
transform 1 0 2632 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_815
timestamp 1543120812
transform 1 0 2520 0 1 870
box -6 -6 6 6
use M3_M2  M3_M2_816
timestamp 1543120812
transform 1 0 2520 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_817
timestamp 1543120812
transform 1 0 2136 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_818
timestamp 1543120812
transform 1 0 1944 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_819
timestamp 1543120812
transform 1 0 1944 0 1 690
box -6 -6 6 6
use M3_M2  M3_M2_820
timestamp 1543120812
transform 1 0 1080 0 1 1210
box -6 -6 6 6
use M3_M2  M3_M2_821
timestamp 1543120812
transform 1 0 1608 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_822
timestamp 1543120812
transform 1 0 1384 0 1 630
box -6 -6 6 6
use M3_M2  M3_M2_823
timestamp 1543120812
transform 1 0 824 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_824
timestamp 1543120812
transform 1 0 600 0 1 1850
box -6 -6 6 6
use M3_M2  M3_M2_825
timestamp 1543120812
transform 1 0 1832 0 1 410
box -6 -6 6 6
use M3_M2  M3_M2_826
timestamp 1543120812
transform 1 0 1528 0 1 410
box -6 -6 6 6
use M3_M2  M3_M2_827
timestamp 1543120812
transform 1 0 1592 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_828
timestamp 1543120812
transform 1 0 1320 0 1 230
box -6 -6 6 6
use M3_M2  M3_M2_829
timestamp 1543120812
transform 1 0 2168 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_830
timestamp 1543120812
transform 1 0 1976 0 1 1990
box -6 -6 6 6
use M3_M2  M3_M2_831
timestamp 1543120812
transform 1 0 1976 0 1 1910
box -6 -6 6 6
use M3_M2  M3_M2_832
timestamp 1543120812
transform 1 0 1384 0 1 1910
box -6 -6 6 6
use M3_M2  M3_M2_833
timestamp 1543120812
transform 1 0 1160 0 1 1910
box -6 -6 6 6
use M3_M2  M3_M2_834
timestamp 1543120812
transform 1 0 1064 0 1 1890
box -6 -6 6 6
use M3_M2  M3_M2_835
timestamp 1543120812
transform 1 0 680 0 1 1890
box -6 -6 6 6
use MUX2X1  MUX2X1_0
timestamp 1053021328
transform 1 0 3408 0 -1 1940
box -10 -6 106 210
use MUX2X1  MUX2X1_1
timestamp 1053021328
transform 1 0 3408 0 1 1540
box -10 -6 106 210
use MUX2X1  MUX2X1_2
timestamp 1053021328
transform 1 0 3264 0 -1 1540
box -10 -6 106 210
use MUX2X1  MUX2X1_3
timestamp 1053021328
transform 1 0 3232 0 1 1140
box -10 -6 106 210
use MUX2X1  MUX2X1_4
timestamp 1053021328
transform 1 0 3472 0 1 1140
box -10 -6 106 210
use MUX2X1  MUX2X1_5
timestamp 1053021328
transform 1 0 3488 0 1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_6
timestamp 1053021328
transform 1 0 3264 0 -1 1140
box -10 -6 106 210
use MUX2X1  MUX2X1_7
timestamp 1053021328
transform 1 0 3264 0 1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_8
timestamp 1053021328
transform 1 0 3248 0 -1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_9
timestamp 1053021328
transform 1 0 3424 0 1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_10
timestamp 1053021328
transform 1 0 3248 0 1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_11
timestamp 1053021328
transform 1 0 3136 0 -1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_12
timestamp 1053021328
transform 1 0 2816 0 1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_13
timestamp 1053021328
transform 1 0 2624 0 -1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_14
timestamp 1053021328
transform 1 0 2848 0 -1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_15
timestamp 1053021328
transform 1 0 2768 0 -1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_16
timestamp 1053021328
transform 1 0 2544 0 -1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_17
timestamp 1053021328
transform 1 0 2272 0 1 340
box -10 -6 106 210
use MUX2X1  MUX2X1_18
timestamp 1053021328
transform 1 0 2320 0 -1 740
box -10 -6 106 210
use MUX2X1  MUX2X1_19
timestamp 1053021328
transform 1 0 2608 0 1 740
box -10 -6 106 210
use NAND2X1  NAND2X1_0
timestamp 1053022145
transform 1 0 2832 0 1 1140
box -16 -6 64 210
use NAND2X1  NAND2X1_1
timestamp 1053022145
transform 1 0 1312 0 -1 1140
box -16 -6 64 210
use NAND2X1  NAND2X1_2
timestamp 1053022145
transform 1 0 1536 0 1 1140
box -16 -6 64 210
use NAND2X1  NAND2X1_3
timestamp 1053022145
transform 1 0 1568 0 1 740
box -16 -6 64 210
use NAND2X1  NAND2X1_4
timestamp 1053022145
transform 1 0 2064 0 1 740
box -16 -6 64 210
use NAND2X1  NAND2X1_5
timestamp 1053022145
transform 1 0 1008 0 -1 1540
box -16 -6 64 210
use NAND2X1  NAND2X1_6
timestamp 1053022145
transform 1 0 592 0 -1 1940
box -16 -6 64 210
use NAND2X1  NAND2X1_7
timestamp 1053022145
transform 1 0 592 0 1 1540
box -16 -6 64 210
use NAND2X1  NAND2X1_8
timestamp 1053022145
transform 1 0 2096 0 1 1140
box -16 -6 64 210
use NAND2X1  NAND2X1_9
timestamp 1053022145
transform 1 0 864 0 1 1540
box -16 -6 64 210
use NAND2X1  NAND2X1_10
timestamp 1053022145
transform 1 0 624 0 1 740
box -16 -6 64 210
use NAND2X1  NAND2X1_11
timestamp 1053022145
transform 1 0 1376 0 -1 740
box -16 -6 64 210
use NAND2X1  NAND2X1_12
timestamp 1053022145
transform 1 0 1424 0 -1 1540
box -16 -6 64 210
use NAND2X1  NAND2X1_13
timestamp 1053022145
transform 1 0 1968 0 -1 1540
box -16 -6 64 210
use NAND2X1  NAND2X1_14
timestamp 1053022145
transform 1 0 1760 0 -1 3540
box -16 -6 64 210
use NAND2X1  NAND2X1_15
timestamp 1053022145
transform 1 0 1632 0 1 2740
box -16 -6 64 210
use NAND2X1  NAND2X1_16
timestamp 1053022145
transform 1 0 2144 0 1 2740
box -16 -6 64 210
use NAND2X1  NAND2X1_17
timestamp 1053022145
transform 1 0 1472 0 1 2740
box -16 -6 64 210
use NAND2X1  NAND2X1_18
timestamp 1053022145
transform 1 0 1872 0 1 2740
box -16 -6 64 210
use NAND2X1  NAND2X1_19
timestamp 1053022145
transform 1 0 1840 0 -1 3140
box -16 -6 64 210
use NAND2X1  NAND2X1_20
timestamp 1053022145
transform 1 0 2208 0 -1 3140
box -16 -6 64 210
use NAND2X1  NAND2X1_21
timestamp 1053022145
transform 1 0 1568 0 -1 3140
box -16 -6 64 210
use NAND2X1  NAND2X1_22
timestamp 1053022145
transform 1 0 2656 0 -1 3140
box -16 -6 64 210
use NAND2X1  NAND2X1_23
timestamp 1053022145
transform 1 0 576 0 -1 3140
box -16 -6 64 210
use NAND3X1  NAND3X1_0
timestamp 1053022145
transform 1 0 448 0 1 740
box -16 -6 80 210
use NAND3X1  NAND3X1_1
timestamp 1053022145
transform 1 0 1104 0 -1 740
box -16 -6 80 210
use NAND3X1  NAND3X1_2
timestamp 1053022145
transform 1 0 880 0 -1 740
box -16 -6 80 210
use NAND3X1  NAND3X1_3
timestamp 1053022145
transform 1 0 1072 0 1 740
box -16 -6 80 210
use NAND3X1  NAND3X1_4
timestamp 1053022145
transform 1 0 928 0 1 1140
box -16 -6 80 210
use NAND3X1  NAND3X1_5
timestamp 1053022145
transform 1 0 1440 0 -1 1140
box -16 -6 80 210
use NAND3X1  NAND3X1_6
timestamp 1053022145
transform 1 0 1744 0 -1 1540
box -16 -6 80 210
use NAND3X1  NAND3X1_7
timestamp 1053022145
transform 1 0 1584 0 -1 3540
box -16 -6 80 210
use NAND3X1  NAND3X1_8
timestamp 1053022145
transform 1 0 400 0 -1 3140
box -16 -6 80 210
use NAND3X1  NAND3X1_9
timestamp 1053022145
transform 1 0 1056 0 -1 3140
box -16 -6 80 210
use NAND3X1  NAND3X1_10
timestamp 1053022145
transform 1 0 992 0 -1 2340
box -16 -6 80 210
use NAND3X1  NAND3X1_11
timestamp 1053022145
transform 1 0 1472 0 1 3140
box -16 -6 80 210
use NAND3X1  NAND3X1_12
timestamp 1053022145
transform 1 0 1008 0 -1 2740
box -16 -6 80 210
use NAND3X1  NAND3X1_13
timestamp 1053022145
transform 1 0 1456 0 -1 340
box -16 -6 80 210
use NOR2X1  NOR2X1_0
timestamp 1053022145
transform 1 0 2496 0 1 340
box -16 -6 64 210
use NOR2X1  NOR2X1_1
timestamp 1053022145
transform 1 0 3024 0 -1 340
box -16 -6 64 210
use NOR2X1  NOR2X1_2
timestamp 1053022145
transform 1 0 3456 0 -1 740
box -16 -6 64 210
use NOR2X1  NOR2X1_3
timestamp 1053022145
transform 1 0 3456 0 -1 1140
box -16 -6 64 210
use NOR2X1  NOR2X1_4
timestamp 1053022145
transform 1 0 3232 0 1 1540
box -16 -6 64 210
use NOR2X1  NOR2X1_5
timestamp 1053022145
transform 1 0 3248 0 -1 1940
box -16 -6 64 210
use NOR2X1  NOR2X1_6
timestamp 1053022145
transform 1 0 512 0 -1 740
box -16 -6 64 210
use NOR2X1  NOR2X1_7
timestamp 1053022145
transform 1 0 512 0 1 740
box -16 -6 64 210
use NOR2X1  NOR2X1_8
timestamp 1053022145
transform 1 0 896 0 -1 1140
box -16 -6 64 210
use NOR2X1  NOR2X1_9
timestamp 1053022145
transform 1 0 1072 0 1 1140
box -16 -6 64 210
use NOR2X1  NOR2X1_10
timestamp 1053022145
transform 1 0 944 0 -1 740
box -16 -6 64 210
use NOR2X1  NOR2X1_11
timestamp 1053022145
transform 1 0 592 0 -1 1540
box -16 -6 64 210
use NOR2X1  NOR2X1_12
timestamp 1053022145
transform 1 0 960 0 -1 1140
box -16 -6 64 210
use NOR2X1  NOR2X1_13
timestamp 1053022145
transform 1 0 1984 0 -1 1140
box -16 -6 64 210
use NOR2X1  NOR2X1_14
timestamp 1053022145
transform 1 0 2544 0 -1 1540
box -16 -6 64 210
use NOR2X1  NOR2X1_15
timestamp 1053022145
transform 1 0 2752 0 1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_16
timestamp 1053022145
transform 1 0 1184 0 1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_17
timestamp 1053022145
transform 1 0 2512 0 1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_18
timestamp 1053022145
transform 1 0 1536 0 -1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_19
timestamp 1053022145
transform 1 0 2480 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_20
timestamp 1053022145
transform 1 0 1184 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_21
timestamp 1053022145
transform 1 0 1936 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_22
timestamp 1053022145
transform 1 0 1344 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_23
timestamp 1053022145
transform 1 0 2320 0 -1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_24
timestamp 1053022145
transform 1 0 1888 0 1 1940
box -16 -6 64 210
use NOR2X1  NOR2X1_25
timestamp 1053022145
transform 1 0 2224 0 1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_26
timestamp 1053022145
transform 1 0 1440 0 1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_27
timestamp 1053022145
transform 1 0 2720 0 1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_28
timestamp 1053022145
transform 1 0 1856 0 -1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_29
timestamp 1053022145
transform 1 0 2752 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_30
timestamp 1053022145
transform 1 0 1664 0 1 2340
box -16 -6 64 210
use NOR2X1  NOR2X1_31
timestamp 1053022145
transform 1 0 2480 0 -1 3140
box -16 -6 64 210
use NOR2X1  NOR2X1_32
timestamp 1053022145
transform 1 0 2496 0 1 1940
box -16 -6 64 210
use NOR2X1  NOR2X1_33
timestamp 1053022145
transform 1 0 2368 0 1 3140
box -16 -6 64 210
use NOR2X1  NOR2X1_34
timestamp 1053022145
transform 1 0 2208 0 -1 2740
box -16 -6 64 210
use NOR2X1  NOR2X1_35
timestamp 1053022145
transform 1 0 1552 0 -1 340
box -16 -6 64 210
use OAI21X1  OAI21X1_0
timestamp 1053722159
transform 1 0 2656 0 1 340
box -16 -6 68 210
use OAI21X1  OAI21X1_1
timestamp 1053722159
transform 1 0 3104 0 1 340
box -16 -6 68 210
use OAI21X1  OAI21X1_2
timestamp 1053722159
transform 1 0 3504 0 -1 740
box -16 -6 68 210
use OAI21X1  OAI21X1_3
timestamp 1053722159
transform 1 0 3360 0 1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_4
timestamp 1053722159
transform 1 0 1248 0 -1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_5
timestamp 1053722159
transform 1 0 1056 0 -1 1540
box -16 -6 68 210
use OAI21X1  OAI21X1_6
timestamp 1053722159
transform 1 0 640 0 1 1540
box -16 -6 68 210
use OAI21X1  OAI21X1_7
timestamp 1053722159
transform 1 0 512 0 -1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_8
timestamp 1053722159
transform 1 0 1168 0 -1 740
box -16 -6 68 210
use OAI21X1  OAI21X1_9
timestamp 1053722159
transform 1 0 672 0 -1 740
box -16 -6 68 210
use OAI21X1  OAI21X1_10
timestamp 1053722159
transform 1 0 736 0 -1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_11
timestamp 1053722159
transform 1 0 672 0 -1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_12
timestamp 1053722159
transform 1 0 816 0 1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_13
timestamp 1053722159
transform 1 0 1136 0 -1 1140
box -16 -6 68 210
use OAI21X1  OAI21X1_14
timestamp 1053722159
transform 1 0 1392 0 1 740
box -16 -6 68 210
use OAI21X1  OAI21X1_15
timestamp 1053722159
transform 1 0 960 0 1 1540
box -16 -6 68 210
use OAI21X1  OAI21X1_16
timestamp 1053722159
transform 1 0 1232 0 -1 1540
box -16 -6 68 210
use OAI21X1  OAI21X1_17
timestamp 1053722159
transform 1 0 1728 0 1 2740
box -16 -6 68 210
use OAI21X1  OAI21X1_18
timestamp 1053722159
transform 1 0 1808 0 1 2740
box -16 -6 68 210
use OAI21X1  OAI21X1_19
timestamp 1053722159
transform 1 0 1968 0 -1 3140
box -16 -6 68 210
use OAI21X1  OAI21X1_20
timestamp 1053722159
transform 1 0 1888 0 -1 3140
box -16 -6 68 210
use OAI22X1  OAI22X1_0
timestamp 1053021427
transform 1 0 1552 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_1
timestamp 1053021427
transform 1 0 1280 0 -1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_2
timestamp 1053021427
transform 1 0 1984 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_3
timestamp 1053021427
transform 1 0 2016 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_4
timestamp 1053021427
transform 1 0 1184 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_5
timestamp 1053021427
transform 1 0 1472 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_6
timestamp 1053021427
transform 1 0 2208 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_7
timestamp 1053021427
transform 1 0 2208 0 -1 1140
box -16 -6 92 210
use OAI22X1  OAI22X1_8
timestamp 1053021427
transform 1 0 1696 0 -1 1140
box -16 -6 92 210
use OAI22X1  OAI22X1_9
timestamp 1053021427
transform 1 0 1696 0 1 1140
box -16 -6 92 210
use OAI22X1  OAI22X1_10
timestamp 1053021427
transform 1 0 1712 0 -1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_11
timestamp 1053021427
transform 1 0 1712 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_12
timestamp 1053021427
transform 1 0 2416 0 -1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_13
timestamp 1053021427
transform 1 0 2464 0 1 1540
box -16 -6 92 210
use OAI22X1  OAI22X1_14
timestamp 1053021427
transform 1 0 2208 0 1 1140
box -16 -6 92 210
use OAI22X1  OAI22X1_15
timestamp 1053021427
transform 1 0 2944 0 -1 2340
box -16 -6 92 210
use OAI22X1  OAI22X1_16
timestamp 1053021427
transform 1 0 864 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_17
timestamp 1053021427
transform 1 0 672 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_18
timestamp 1053021427
transform 1 0 2928 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_19
timestamp 1053021427
transform 1 0 3024 0 1 2740
box -16 -6 92 210
use OAI22X1  OAI22X1_20
timestamp 1053021427
transform 1 0 1136 0 -1 3540
box -16 -6 92 210
use OAI22X1  OAI22X1_21
timestamp 1053021427
transform 1 0 752 0 -1 3140
box -16 -6 92 210
use OAI22X1  OAI22X1_22
timestamp 1053021427
transform 1 0 3168 0 -1 3140
box -16 -6 92 210
use OAI22X1  OAI22X1_23
timestamp 1053021427
transform 1 0 2480 0 -1 3540
box -16 -6 92 210
use OAI22X1  OAI22X1_24
timestamp 1053021427
transform 1 0 3072 0 -1 3540
box -16 -6 92 210
use OAI22X1  OAI22X1_25
timestamp 1053021427
transform 1 0 2784 0 -1 3540
box -16 -6 92 210
use OAI22X1  OAI22X1_26
timestamp 1053021427
transform 1 0 2112 0 -1 3540
box -16 -6 92 210
use OAI22X1  OAI22X1_27
timestamp 1053021427
transform 1 0 3248 0 1 2740
box -16 -6 92 210
use OAI22X1  OAI22X1_28
timestamp 1053021427
transform 1 0 672 0 1 2340
box -16 -6 92 210
use OAI22X1  OAI22X1_29
timestamp 1053021427
transform 1 0 592 0 -1 2740
box -16 -6 92 210
use OAI22X1  OAI22X1_30
timestamp 1053021427
transform 1 0 2992 0 1 2340
box -16 -6 92 210
use OAI22X1  OAI22X1_31
timestamp 1053021427
transform 1 0 2064 0 1 1940
box -16 -6 92 210
use OAI22X1  OAI22X1_32
timestamp 1053021427
transform 1 0 752 0 1 3140
box -16 -6 92 210
use OR2X1  OR2X1_0
timestamp 1090542464
transform 1 0 2896 0 1 740
box -16 -6 80 210
use OR2X1  OR2X1_1
timestamp 1090542464
transform 1 0 3088 0 1 1540
box -16 -6 80 210
use OR2X1  OR2X1_2
timestamp 1090542464
transform 1 0 3024 0 1 1540
box -16 -6 80 210
use OR2X1  OR2X1_3
timestamp 1090542464
transform 1 0 3104 0 1 1140
box -16 -6 80 210
use OR2X1  OR2X1_4
timestamp 1090542464
transform 1 0 3136 0 -1 1140
box -16 -6 80 210
use OR2X1  OR2X1_5
timestamp 1090542464
transform 1 0 3152 0 1 740
box -16 -6 80 210
use OR2X1  OR2X1_6
timestamp 1090542464
transform 1 0 2864 0 -1 740
box -16 -6 80 210
use OR2X1  OR2X1_7
timestamp 1090542464
transform 1 0 672 0 1 1140
box -16 -6 80 210
use top_VIA0  top_VIA0_0
timestamp 1543120812
transform 1 0 3776 0 1 3634
box -20 -20 20 20
use top_VIA0  top_VIA0_1
timestamp 1543120812
transform 1 0 3776 0 1 46
box -20 -20 20 20
use top_VIA0  top_VIA0_2
timestamp 1543120812
transform 1 0 48 0 1 3634
box -20 -20 20 20
use top_VIA0  top_VIA0_3
timestamp 1543120812
transform 1 0 48 0 1 46
box -20 -20 20 20
use top_VIA0  top_VIA0_4
timestamp 1543120812
transform 1 0 3728 0 1 3586
box -20 -20 20 20
use top_VIA0  top_VIA0_5
timestamp 1543120812
transform 1 0 3728 0 1 94
box -20 -20 20 20
use top_VIA0  top_VIA0_6
timestamp 1543120812
transform 1 0 96 0 1 3586
box -20 -20 20 20
use top_VIA0  top_VIA0_7
timestamp 1543120812
transform 1 0 96 0 1 94
box -20 -20 20 20
use top_VIA1  top_VIA1_0
timestamp 1543120812
transform 1 0 3776 0 1 3340
box -20 -6 20 6
use top_VIA1  top_VIA1_1
timestamp 1543120812
transform 1 0 3776 0 1 2940
box -20 -6 20 6
use top_VIA1  top_VIA1_2
timestamp 1543120812
transform 1 0 3776 0 1 2540
box -20 -6 20 6
use top_VIA1  top_VIA1_3
timestamp 1543120812
transform 1 0 3776 0 1 2140
box -20 -6 20 6
use top_VIA1  top_VIA1_4
timestamp 1543120812
transform 1 0 3776 0 1 1740
box -20 -6 20 6
use top_VIA1  top_VIA1_5
timestamp 1543120812
transform 1 0 3776 0 1 1340
box -20 -6 20 6
use top_VIA1  top_VIA1_6
timestamp 1543120812
transform 1 0 3776 0 1 940
box -20 -6 20 6
use top_VIA1  top_VIA1_7
timestamp 1543120812
transform 1 0 3776 0 1 540
box -20 -6 20 6
use top_VIA1  top_VIA1_8
timestamp 1543120812
transform 1 0 3776 0 1 140
box -20 -6 20 6
use top_VIA1  top_VIA1_9
timestamp 1543120812
transform 1 0 48 0 1 3340
box -20 -6 20 6
use top_VIA1  top_VIA1_10
timestamp 1543120812
transform 1 0 48 0 1 2940
box -20 -6 20 6
use top_VIA1  top_VIA1_11
timestamp 1543120812
transform 1 0 48 0 1 2540
box -20 -6 20 6
use top_VIA1  top_VIA1_12
timestamp 1543120812
transform 1 0 48 0 1 2140
box -20 -6 20 6
use top_VIA1  top_VIA1_13
timestamp 1543120812
transform 1 0 48 0 1 1740
box -20 -6 20 6
use top_VIA1  top_VIA1_14
timestamp 1543120812
transform 1 0 48 0 1 1340
box -20 -6 20 6
use top_VIA1  top_VIA1_15
timestamp 1543120812
transform 1 0 48 0 1 940
box -20 -6 20 6
use top_VIA1  top_VIA1_16
timestamp 1543120812
transform 1 0 48 0 1 540
box -20 -6 20 6
use top_VIA1  top_VIA1_17
timestamp 1543120812
transform 1 0 48 0 1 140
box -20 -6 20 6
use top_VIA1  top_VIA1_18
timestamp 1543120812
transform 1 0 96 0 1 340
box -20 -6 20 6
use top_VIA1  top_VIA1_19
timestamp 1543120812
transform 1 0 96 0 1 740
box -20 -6 20 6
use top_VIA1  top_VIA1_20
timestamp 1543120812
transform 1 0 96 0 1 1140
box -20 -6 20 6
use top_VIA1  top_VIA1_21
timestamp 1543120812
transform 1 0 96 0 1 1540
box -20 -6 20 6
use top_VIA1  top_VIA1_22
timestamp 1543120812
transform 1 0 96 0 1 1940
box -20 -6 20 6
use top_VIA1  top_VIA1_23
timestamp 1543120812
transform 1 0 96 0 1 2340
box -20 -6 20 6
use top_VIA1  top_VIA1_24
timestamp 1543120812
transform 1 0 96 0 1 2740
box -20 -6 20 6
use top_VIA1  top_VIA1_25
timestamp 1543120812
transform 1 0 96 0 1 3140
box -20 -6 20 6
use top_VIA1  top_VIA1_26
timestamp 1543120812
transform 1 0 96 0 1 3540
box -20 -6 20 6
use top_VIA1  top_VIA1_27
timestamp 1543120812
transform 1 0 3728 0 1 340
box -20 -6 20 6
use top_VIA1  top_VIA1_28
timestamp 1543120812
transform 1 0 3728 0 1 740
box -20 -6 20 6
use top_VIA1  top_VIA1_29
timestamp 1543120812
transform 1 0 3728 0 1 1140
box -20 -6 20 6
use top_VIA1  top_VIA1_30
timestamp 1543120812
transform 1 0 3728 0 1 1540
box -20 -6 20 6
use top_VIA1  top_VIA1_31
timestamp 1543120812
transform 1 0 3728 0 1 1940
box -20 -6 20 6
use top_VIA1  top_VIA1_32
timestamp 1543120812
transform 1 0 3728 0 1 2340
box -20 -6 20 6
use top_VIA1  top_VIA1_33
timestamp 1543120812
transform 1 0 3728 0 1 2740
box -20 -6 20 6
use top_VIA1  top_VIA1_34
timestamp 1543120812
transform 1 0 3728 0 1 3140
box -20 -6 20 6
use top_VIA1  top_VIA1_35
timestamp 1543120812
transform 1 0 3728 0 1 3540
box -20 -6 20 6
use XNOR2X1  XNOR2X1_0
timestamp 1054159935
transform 1 0 2368 0 1 340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_1
timestamp 1054159935
transform 1 0 2640 0 -1 740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_2
timestamp 1054159935
transform 1 0 2720 0 -1 340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_3
timestamp 1054159935
transform 1 0 2912 0 1 340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_4
timestamp 1054159935
transform 1 0 3520 0 1 340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_5
timestamp 1054159935
transform 1 0 3344 0 -1 740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_6
timestamp 1054159935
transform 1 0 3504 0 -1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_7
timestamp 1054159935
transform 1 0 3568 0 1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_8
timestamp 1054159935
transform 1 0 3296 0 1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_9
timestamp 1054159935
transform 1 0 3296 0 -1 1940
box -16 -6 128 210
use XNOR2X1  XNOR2X1_10
timestamp 1054159935
transform 1 0 2992 0 1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_11
timestamp 1054159935
transform 1 0 1984 0 1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_12
timestamp 1054159935
transform 1 0 2032 0 -1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_13
timestamp 1054159935
transform 1 0 1504 0 -1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_14
timestamp 1054159935
transform 1 0 1424 0 1 1140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_15
timestamp 1054159935
transform 1 0 2592 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_16
timestamp 1054159935
transform 1 0 2432 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_17
timestamp 1054159935
transform 1 0 1808 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_18
timestamp 1054159935
transform 1 0 1600 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_19
timestamp 1054159935
transform 1 0 1312 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_20
timestamp 1054159935
transform 1 0 1472 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_21
timestamp 1054159935
transform 1 0 2016 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_22
timestamp 1054159935
transform 1 0 2128 0 -1 1540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_23
timestamp 1054159935
transform 1 0 1648 0 -1 3540
box -16 -6 128 210
use XNOR2X1  XNOR2X1_24
timestamp 1054159935
transform 1 0 2528 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_25
timestamp 1054159935
transform 1 0 2640 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_26
timestamp 1054159935
transform 1 0 1072 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_27
timestamp 1054159935
transform 1 0 960 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_28
timestamp 1054159935
transform 1 0 2560 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_29
timestamp 1054159935
transform 1 0 2400 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_30
timestamp 1054159935
transform 1 0 1424 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_31
timestamp 1054159935
transform 1 0 1296 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_32
timestamp 1054159935
transform 1 0 1248 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_33
timestamp 1054159935
transform 1 0 1520 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_34
timestamp 1054159935
transform 1 0 2032 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_35
timestamp 1054159935
transform 1 0 2192 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_36
timestamp 1054159935
transform 1 0 2528 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_37
timestamp 1054159935
transform 1 0 2416 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_38
timestamp 1054159935
transform 1 0 1072 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_39
timestamp 1054159935
transform 1 0 848 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_40
timestamp 1054159935
transform 1 0 2368 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_41
timestamp 1054159935
transform 1 0 1984 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_42
timestamp 1054159935
transform 1 0 1200 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_43
timestamp 1054159935
transform 1 0 1232 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_44
timestamp 1054159935
transform 1 0 1360 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_45
timestamp 1054159935
transform 1 0 1392 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_46
timestamp 1054159935
transform 1 0 1920 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_47
timestamp 1054159935
transform 1 0 2304 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_48
timestamp 1054159935
transform 1 0 2512 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_49
timestamp 1054159935
transform 1 0 2368 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_50
timestamp 1054159935
transform 1 0 1664 0 1 1940
box -16 -6 128 210
use XNOR2X1  XNOR2X1_51
timestamp 1054159935
transform 1 0 1776 0 1 1940
box -16 -6 128 210
use XNOR2X1  XNOR2X1_52
timestamp 1054159935
transform 1 0 2272 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_53
timestamp 1054159935
transform 1 0 2112 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_54
timestamp 1054159935
transform 1 0 1328 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_55
timestamp 1054159935
transform 1 0 1504 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_56
timestamp 1054159935
transform 1 0 1616 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_57
timestamp 1054159935
transform 1 0 1728 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_58
timestamp 1054159935
transform 1 0 2096 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_59
timestamp 1054159935
transform 1 0 2256 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_60
timestamp 1054159935
transform 1 0 2768 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_61
timestamp 1054159935
transform 1 0 2704 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_62
timestamp 1054159935
transform 1 0 1632 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_63
timestamp 1054159935
transform 1 0 1744 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_64
timestamp 1054159935
transform 1 0 2800 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_65
timestamp 1054159935
transform 1 0 2640 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_66
timestamp 1054159935
transform 1 0 1552 0 1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_67
timestamp 1054159935
transform 1 0 1616 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_68
timestamp 1054159935
transform 1 0 1344 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_69
timestamp 1054159935
transform 1 0 1456 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_70
timestamp 1054159935
transform 1 0 2704 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_71
timestamp 1054159935
transform 1 0 2816 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_72
timestamp 1054159935
transform 1 0 464 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_73
timestamp 1054159935
transform 1 0 544 0 1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_74
timestamp 1054159935
transform 1 0 544 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_75
timestamp 1054159935
transform 1 0 864 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_76
timestamp 1054159935
transform 1 0 2528 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_77
timestamp 1054159935
transform 1 0 2368 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_78
timestamp 1054159935
transform 1 0 1120 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_79
timestamp 1054159935
transform 1 0 1232 0 -1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_80
timestamp 1054159935
transform 1 0 2544 0 1 1940
box -16 -6 128 210
use XNOR2X1  XNOR2X1_81
timestamp 1054159935
transform 1 0 2384 0 1 1940
box -16 -6 128 210
use XNOR2X1  XNOR2X1_82
timestamp 1054159935
transform 1 0 880 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_83
timestamp 1054159935
transform 1 0 1104 0 -1 2340
box -16 -6 128 210
use XNOR2X1  XNOR2X1_84
timestamp 1054159935
transform 1 0 2640 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_85
timestamp 1054159935
transform 1 0 2256 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_86
timestamp 1054159935
transform 1 0 1360 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_87
timestamp 1054159935
transform 1 0 1536 0 1 3140
box -16 -6 128 210
use XNOR2X1  XNOR2X1_88
timestamp 1054159935
transform 1 0 2256 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_89
timestamp 1054159935
transform 1 0 2096 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_90
timestamp 1054159935
transform 1 0 896 0 -1 2740
box -16 -6 128 210
use XNOR2X1  XNOR2X1_91
timestamp 1054159935
transform 1 0 1040 0 1 2340
box -16 -6 128 210
use XOR2X1  XOR2X1_0
timestamp 1053359338
transform 1 0 2880 0 1 1140
box -16 -6 128 210
use XOR2X1  XOR2X1_1
timestamp 1053359338
transform 1 0 2928 0 -1 1540
box -16 -6 128 210
use XOR2X1  XOR2X1_2
timestamp 1053359338
transform 1 0 1840 0 -1 3540
box -16 -6 128 210
use XOR2X1  XOR2X1_3
timestamp 1053359338
transform 1 0 1728 0 1 3140
box -16 -6 128 210
use XOR2X1  XOR2X1_4
timestamp 1053359338
transform 1 0 1920 0 1 3140
box -16 -6 128 210
<< labels >>
rlabel metal1 2232 1870 2232 1870 4 in_clka
rlabel electrodecontact s 3256 1990 3256 1990 4 in_clkb
rlabel electrodecontact s 1496 210 1496 210 4 in_enter
rlabel metal1 1752 270 1752 270 4 in_restart
rlabel electrodecontact s 2200 3470 2200 3470 4 in_ans0[3]
rlabel electrodecontact s 2872 3470 2872 3470 4 in_ans0[2]
rlabel electrodecontact s 3224 3470 3224 3470 4 in_ans0[1]
rlabel electrodecontact s 2456 3470 2456 3470 4 in_ans0[0]
rlabel electrodecontact s 3288 3070 3288 3070 4 in_ans1[3]
rlabel electrodecontact s 728 3070 728 3070 4 in_ans1[2]
rlabel electrodecontact s 1224 3470 1224 3470 4 in_ans1[1]
rlabel electrodecontact s 3112 2810 3112 2810 4 in_ans1[0]
rlabel electrodecontact s 3048 2010 3048 2010 4 in_ans2[3]
rlabel electrodecontact s 648 2010 648 2010 4 in_ans2[2]
rlabel electrodecontact s 840 2010 840 2010 4 in_ans2[1]
rlabel electrodecontact s 2920 2270 2920 2270 4 in_ans2[0]
rlabel electrodecontact s 3080 2410 3080 2410 4 in_ans3[3]
rlabel electrodecontact s 536 2670 536 2670 4 in_ans3[2]
rlabel electrodecontact s 584 2410 584 2410 4 in_ans3[1]
rlabel electrodecontact s 3352 2810 3352 2810 4 in_ans3[0]
rlabel electrodecontact s 376 3050 376 3050 4 out_Anum[2]
rlabel electrodecontact s 536 3050 536 3050 4 out_Anum[1]
rlabel electrodecontact s 616 2830 616 2830 4 out_Anum[0]
rlabel electrodecontact s 1496 3450 1496 3450 4 out_Bnum[2]
rlabel electrodecontact s 1720 3450 1720 3450 4 out_Bnum[1]
rlabel electrodecontact s 1896 3450 1896 3450 4 out_Bnum[0]
rlabel electrodecontact s 1320 250 1320 250 4 out_state[1]
rlabel metal1 1624 410 1624 410 4 out_state[0]
rlabel electrodecontact s 840 1850 840 1850 4 out_valid
rlabel metal2 76 74 76 74 4 gnd
rlabel metal2 28 26 28 26 4 vdd
<< properties >>
string path 6102.000 922.500 6180.750 922.500 
<< end >>
