* SPICE3 file created from top.ext - technology: scmos

.option scale=0.3u

M1000 DFFNEGX1_40/a_76_6# INVX4_0/Y DFFNEGX1_40/a_66_6# Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=40p ps=18u
M1001 gnd INVX4_0/Y DFFNEGX1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=55p pd=26u as=100p ps=50u
M1002 DFFNEGX1_40/a_66_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_61_6# Gnd nfet w=10 l=2
+  ad=40p pd=18u as=14.999999p ps=13u
M1003 INVX2_57/A DFFNEGX1_40/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=55p ps=26u
M1004 DFFNEGX1_40/a_23_6# INVX4_0/Y DFFNEGX1_40/a_17_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=20p ps=14u
M1005 DFFNEGX1_40/a_23_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_17_74# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=40p ps=24u
M1006 gnd DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_31_6# Gnd nfet w=10 l=2
+  ad=35p pd=17u as=14.999999p ps=13u
M1007 vdd DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_31_74# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=40p ps=24u
M1008 DFFNEGX1_40/a_61_74# DFFNEGX1_40/a_34_4# vdd vdd pfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1009 DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1010 DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=35p ps=17u
M1011 vdd INVX2_57/A DFFNEGX1_40/a_76_84# vdd pfet w=10 l=2
+  ad=0.105n pd=46u as=14.999999p ps=13u
M1012 gnd INVX2_57/A DFFNEGX1_40/a_76_6# Gnd nfet w=10 l=2
+  ad=55p pd=26u as=14.999999p ps=13u
M1013 DFFNEGX1_40/a_61_6# DFFNEGX1_40/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=50p ps=30u
M1014 DFFNEGX1_40/a_76_84# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_66_6# vdd pfet w=10 l=2
+  ad=14.999999p pd=13u as=75p ps=28u
M1015 INVX2_57/A DFFNEGX1_40/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.105n ps=46u
M1016 vdd INVX4_0/Y DFFNEGX1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=0.2n ps=90u
M1017 DFFNEGX1_40/a_31_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_23_6# Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=29.999998p ps=16u
M1018 DFFNEGX1_40/a_66_6# INVX4_0/Y DFFNEGX1_40/a_61_74# vdd pfet w=20 l=2
+  ad=75p pd=28u as=29.999998p ps=23u
M1019 DFFNEGX1_40/a_17_74# OAI22X1_23/Y vdd vdd pfet w=20 l=2
+  ad=40p pd=24u as=0.11n ps=46u
M1020 DFFNEGX1_40/a_31_74# INVX4_0/Y DFFNEGX1_40/a_23_6# vdd pfet w=20 l=2
+  ad=40p pd=24u as=59.999996p ps=26u
M1021 DFFNEGX1_40/a_17_6# OAI22X1_23/Y gnd Gnd nfet w=10 l=2
+  ad=20p pd=14u as=55p ps=26u
M1022 gnd XNOR2X1_0/Y MUX2X1_17/a_30_10# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1023 MUX2X1_17/a_17_50# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.104n ps=46u
M1024 INVX2_15/A OAI21X1_0/Y MUX2X1_17/a_17_50# vdd pfet w=40 l=2
+  ad=0.124n pd=50u as=59.999996p ps=43u
M1025 MUX2X1_17/a_30_54# MUX2X1_17/a_2_10# INVX2_15/A vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.124n ps=50u
M1026 MUX2X1_17/a_17_10# NOR2X1_0/A gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=53p ps=26u
M1027 vdd OAI21X1_0/Y MUX2X1_17/a_2_10# vdd pfet w=20 l=2
+  ad=0.104n pd=46u as=100p ps=50u
M1028 MUX2X1_17/a_30_10# OAI21X1_0/Y INVX2_15/A Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=59.999996p ps=26u
M1029 gnd OAI21X1_0/Y MUX2X1_17/a_2_10# Gnd nfet w=10 l=2
+  ad=53p pd=26u as=50p ps=30u
M1030 vdd XNOR2X1_0/Y MUX2X1_17/a_30_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M1031 INVX2_15/A MUX2X1_17/a_2_10# MUX2X1_17/a_17_10# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=29.999998p ps=23u
M1032 gnd NAND2X1_4/A AOI22X1_0/a_28_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1033 INVX2_74/A DFFSR_7/S AOI22X1_0/a_11_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M1034 AOI22X1_0/a_11_6# INVX2_14/Y gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1035 AOI22X1_0/a_2_54# DFFSR_7/S vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1036 AOI22X1_0/a_28_6# INVX2_99/A INVX2_74/A Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M1037 vdd INVX2_14/Y AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M1038 INVX2_74/A INVX2_99/A AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1039 AOI22X1_0/a_2_54# NAND2X1_4/A INVX2_74/A vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M1040 OAI21X1_14/A XNOR2X1_13/Y vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1041 NAND2X1_10/a_9_6# XNOR2X1_13/Y gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1042 vdd XNOR2X1_12/Y OAI21X1_14/A vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1043 OAI21X1_14/A XNOR2X1_12/Y NAND2X1_10/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1044 OAI21X1_20/A XNOR2X1_70/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0.16143u ps=0.066482
M1045 NAND2X1_21/a_9_6# XNOR2X1_70/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=79.270004n ps=0.035986
M1046 vdd XNOR2X1_69/Y OAI21X1_20/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1047 OAI21X1_20/A XNOR2X1_69/Y NAND2X1_21/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1048 gnd OAI22X1_6/A OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1049 OAI22X1_3/a_2_6# INVX2_98/Y OAI22X1_3/Y Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1050 OAI22X1_3/Y INVX2_78/Y OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1051 OAI22X1_3/Y INVX2_42/Y OAI22X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0.24n pd=52u as=59.999996p ps=43u
M1052 OAI22X1_3/a_28_54# INVX2_78/Y OAI22X1_3/Y vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.24n ps=52u
M1053 OAI22X1_3/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M1054 OAI22X1_3/a_2_6# INVX2_42/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1055 vdd INVX2_98/Y OAI22X1_3/a_28_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M1056 NOR2X1_0/A INVX2_12/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1057 NOR2X1_0/A INVX2_12/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1058 INVX2_34/Y INVX2_34/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1059 INVX2_34/Y INVX2_34/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1060 INVX2_23/Y INVX2_23/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1061 INVX2_23/Y INVX2_23/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1062 INVX2_67/Y INVX2_67/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1063 INVX2_67/Y INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1064 INVX2_45/Y INVX2_45/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1065 INVX2_45/Y INVX2_45/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1066 INVX2_78/Y in_ans3[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1067 INVX2_78/Y in_ans3[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1068 INVX2_56/Y INVX2_56/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1069 INVX2_56/Y INVX2_56/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1070 INVX2_89/Y in_ans1[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1071 INVX2_89/Y in_ans1[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1072 gnd OAI21X1_19/A OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1073 vdd AOI22X1_7/Y XOR2X1_5/A vdd pfet w=20 l=2
+  ad=100p pd=50u as=0.11n ps=46u
M1074 XOR2X1_5/A AOI22X1_7/Y OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1075 XOR2X1_5/A OAI21X1_19/B OAI21X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=59.999996p ps=43u
M1076 OAI21X1_19/a_9_54# OAI21X1_19/A vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M1077 OAI21X1_19/a_2_6# OAI21X1_19/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1078 gnd INVX2_4/Y XNOR2X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=100p ps=50u
M1079 MUX2X1_5/A INVX2_4/Y XNOR2X1_6/a_18_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M1080 XNOR2X1_6/a_12_41# INVX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=70p ps=27u
M1081 XNOR2X1_6/a_18_54# XNOR2X1_6/a_12_41# vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.14n ps=47u
M1082 XNOR2X1_6/a_35_6# XNOR2X1_6/a_2_6# MUX2X1_5/A Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M1083 XNOR2X1_6/a_18_6# XNOR2X1_6/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=70p ps=27u
M1084 vdd INVX2_4/Y XNOR2X1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=0.2n ps=90u
M1085 vdd INVX2_3/Y XNOR2X1_6/a_35_54# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=59.999996p ps=43u
M1086 MUX2X1_5/A XNOR2X1_6/a_2_6# XNOR2X1_6/a_18_54# vdd pfet w=40 l=2
+  ad=0.2n pd=50u as=59.999996p ps=43u
M1087 XNOR2X1_6/a_35_54# INVX2_4/Y MUX2X1_5/A vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=50u
M1088 XNOR2X1_6/a_12_41# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.14n ps=47u
M1089 gnd INVX2_3/Y XNOR2X1_6/a_35_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=29.999998p ps=23u
M1090 DFFNEGX1_41/a_76_6# INVX2_102/Y DFFNEGX1_41/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1091 gnd INVX2_102/Y DFFNEGX1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1092 DFFNEGX1_41/a_66_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1093 out_state[0] DFFNEGX1_41/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1094 DFFNEGX1_41/a_23_6# INVX2_102/Y DFFNEGX1_41/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1095 DFFNEGX1_41/a_23_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1096 gnd DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1097 vdd DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1098 DFFNEGX1_41/a_61_74# DFFNEGX1_41/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1099 DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1100 DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1101 vdd out_state[0] DFFNEGX1_41/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1102 gnd out_state[0] DFFNEGX1_41/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1103 DFFNEGX1_41/a_61_6# DFFNEGX1_41/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1104 DFFNEGX1_41/a_76_84# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1105 out_state[0] DFFNEGX1_41/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1106 vdd INVX2_102/Y DFFNEGX1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1107 DFFNEGX1_41/a_31_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 DFFNEGX1_41/a_66_6# INVX2_102/Y DFFNEGX1_41/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 DFFNEGX1_41/a_17_74# AND2X2_4/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 DFFNEGX1_41/a_31_74# INVX2_102/Y DFFNEGX1_41/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1111 DFFNEGX1_41/a_17_6# AND2X2_4/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 DFFNEGX1_30/a_76_6# INVX4_0/Y DFFNEGX1_30/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1113 gnd INVX4_0/Y DFFNEGX1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1114 DFFNEGX1_30/a_66_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1115 INVX2_45/A DFFNEGX1_30/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1116 DFFNEGX1_30/a_23_6# INVX4_0/Y DFFNEGX1_30/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1117 DFFNEGX1_30/a_23_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1118 gnd DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1119 vdd DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1120 DFFNEGX1_30/a_61_74# DFFNEGX1_30/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1121 DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1122 DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1123 vdd INVX2_45/A DFFNEGX1_30/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1124 gnd INVX2_45/A DFFNEGX1_30/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1125 DFFNEGX1_30/a_61_6# DFFNEGX1_30/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1126 DFFNEGX1_30/a_76_84# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1127 INVX2_45/A DFFNEGX1_30/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1128 vdd INVX4_0/Y DFFNEGX1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1129 DFFNEGX1_30/a_31_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 DFFNEGX1_30/a_66_6# INVX4_0/Y DFFNEGX1_30/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 DFFNEGX1_30/a_17_74# OAI22X1_1/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 DFFNEGX1_30/a_31_74# INVX4_0/Y DFFNEGX1_30/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 DFFNEGX1_30/a_17_6# OAI22X1_1/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1134 gnd INVX2_13/A MUX2X1_18/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1135 MUX2X1_18/a_17_50# NOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1136 INVX2_16/A OAI21X1_0/Y MUX2X1_18/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1137 MUX2X1_18/a_30_54# MUX2X1_18/a_2_10# INVX2_16/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1138 MUX2X1_18/a_17_10# NOR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1139 vdd OAI21X1_0/Y MUX2X1_18/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1140 MUX2X1_18/a_30_10# OAI21X1_0/Y INVX2_16/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1141 gnd OAI21X1_0/Y MUX2X1_18/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1142 vdd INVX2_13/A MUX2X1_18/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1143 INVX2_16/A MUX2X1_18/a_2_10# MUX2X1_18/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 gnd NAND2X1_3/A AOI22X1_1/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1145 INVX2_75/A DFFSR_7/S AOI22X1_1/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1146 AOI22X1_1/a_11_6# INVX2_15/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 AOI22X1_1/a_2_54# DFFSR_7/S vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1148 AOI22X1_1/a_28_6# INVX2_99/A INVX2_75/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1149 vdd INVX2_15/Y AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1150 INVX2_75/A INVX2_99/A AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1151 AOI22X1_1/a_2_54# NAND2X1_3/A INVX2_75/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 OAI22X1_7/D AOI22X1_3/C vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1153 NAND2X1_11/a_9_6# AOI22X1_3/C gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1154 vdd INVX2_72/Y OAI22X1_7/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1155 OAI22X1_7/D INVX2_72/Y NAND2X1_11/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1156 XNOR2X1_71/A INVX2_43/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1157 NAND2X1_22/a_9_6# INVX2_43/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1158 vdd NAND3X1_8/A XNOR2X1_71/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 XNOR2X1_71/A NAND3X1_8/A NAND2X1_22/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1160 gnd OAI22X1_6/A OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1161 OAI22X1_4/a_2_6# INVX2_98/Y OAI22X1_4/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1162 OAI22X1_4/Y INVX2_79/Y OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1163 OAI22X1_4/Y INVX2_41/Y OAI22X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1164 OAI22X1_4/a_28_54# INVX2_79/Y OAI22X1_4/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1165 OAI22X1_4/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 OAI22X1_4/a_2_6# INVX2_41/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 vdd INVX2_98/Y OAI22X1_4/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1168 NOR2X1_0/B INVX2_13/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1169 NOR2X1_0/B INVX2_13/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1170 INVX2_68/Y INVX2_68/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1171 INVX2_68/Y INVX2_68/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1172 INVX2_24/Y INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1173 INVX2_24/Y INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1174 INVX2_57/Y INVX2_57/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1175 INVX2_57/Y INVX2_57/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1176 INVX2_79/Y in_ans3[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1177 INVX2_79/Y in_ans3[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1178 INVX2_46/Y INVX2_46/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1179 INVX2_46/Y INVX2_46/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1180 INVX2_35/Y INVX2_35/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1181 INVX2_35/Y INVX2_35/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1182 gnd INVX2_2/Y XNOR2X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1183 MUX2X1_4/A INVX2_2/Y XNOR2X1_7/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1184 XNOR2X1_7/a_12_41# NOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1185 XNOR2X1_7/a_18_54# XNOR2X1_7/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1186 XNOR2X1_7/a_35_6# XNOR2X1_7/a_2_6# MUX2X1_4/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1187 XNOR2X1_7/a_18_6# XNOR2X1_7/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 vdd INVX2_2/Y XNOR2X1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1189 vdd NOR2X1_3/Y XNOR2X1_7/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1190 MUX2X1_4/A XNOR2X1_7/a_2_6# XNOR2X1_7/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1191 XNOR2X1_7/a_35_54# INVX2_2/Y MUX2X1_4/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 XNOR2X1_7/a_12_41# NOR2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1193 gnd NOR2X1_3/Y XNOR2X1_7/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 DFFNEGX1_42/a_76_6# in_clka DFFNEGX1_42/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1195 gnd in_clka DFFNEGX1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1196 DFFNEGX1_42/a_66_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1197 out_state[1] DFFNEGX1_42/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1198 DFFNEGX1_42/a_23_6# in_clka DFFNEGX1_42/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1199 DFFNEGX1_42/a_23_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1200 gnd DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1201 vdd DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1202 DFFNEGX1_42/a_61_74# DFFNEGX1_42/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1203 DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1204 DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1205 vdd out_state[1] DFFNEGX1_42/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1206 gnd out_state[1] DFFNEGX1_42/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1207 DFFNEGX1_42/a_61_6# DFFNEGX1_42/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 DFFNEGX1_42/a_76_84# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1209 out_state[1] DFFNEGX1_42/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1210 vdd in_clka DFFNEGX1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1211 DFFNEGX1_42/a_31_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1212 DFFNEGX1_42/a_66_6# in_clka DFFNEGX1_42/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 DFFNEGX1_42/a_17_74# NOR2X1_37/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 DFFNEGX1_42/a_31_74# in_clka DFFNEGX1_42/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 DFFNEGX1_42/a_17_6# NOR2X1_37/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 DFFNEGX1_20/a_76_6# INVX2_102/Y DFFNEGX1_20/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1217 gnd INVX2_102/Y DFFNEGX1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1218 DFFNEGX1_20/a_66_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1219 out_valid DFFNEGX1_20/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1220 DFFNEGX1_20/a_23_6# INVX2_102/Y DFFNEGX1_20/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1221 DFFNEGX1_20/a_23_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1222 gnd DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1223 vdd DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1224 DFFNEGX1_20/a_61_74# DFFNEGX1_20/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1225 DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1226 DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1227 vdd out_valid DFFNEGX1_20/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1228 gnd out_valid DFFNEGX1_20/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1229 DFFNEGX1_20/a_61_6# DFFNEGX1_20/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 DFFNEGX1_20/a_76_84# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1231 out_valid DFFNEGX1_20/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1232 vdd INVX2_102/Y DFFNEGX1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1233 DFFNEGX1_20/a_31_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 DFFNEGX1_20/a_66_6# INVX2_102/Y DFFNEGX1_20/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 DFFNEGX1_20/a_17_74# OAI21X1_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1236 DFFNEGX1_20/a_31_74# INVX2_102/Y DFFNEGX1_20/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1237 DFFNEGX1_20/a_17_6# OAI21X1_7/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1238 DFFNEGX1_31/a_76_6# INVX4_0/Y DFFNEGX1_31/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1239 gnd INVX4_0/Y DFFNEGX1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1240 DFFNEGX1_31/a_66_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1241 INVX2_46/A DFFNEGX1_31/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1242 DFFNEGX1_31/a_23_6# INVX4_0/Y DFFNEGX1_31/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1243 DFFNEGX1_31/a_23_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1244 gnd DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1245 vdd DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1246 DFFNEGX1_31/a_61_74# DFFNEGX1_31/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1247 DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1248 DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1249 vdd INVX2_46/A DFFNEGX1_31/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1250 gnd INVX2_46/A DFFNEGX1_31/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 DFFNEGX1_31/a_61_6# DFFNEGX1_31/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1252 DFFNEGX1_31/a_76_84# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1253 INVX2_46/A DFFNEGX1_31/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1254 vdd INVX4_0/Y DFFNEGX1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1255 DFFNEGX1_31/a_31_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1256 DFFNEGX1_31/a_66_6# INVX4_0/Y DFFNEGX1_31/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1257 DFFNEGX1_31/a_17_74# OAI22X1_0/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1258 DFFNEGX1_31/a_31_74# INVX4_0/Y DFFNEGX1_31/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 DFFNEGX1_31/a_17_6# OAI22X1_0/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1260 gnd DFFSR_1/D MUX2X1_19/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1261 MUX2X1_19/a_17_50# DFFSR_1/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1262 INVX2_17/A OAI21X1_0/Y MUX2X1_19/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1263 MUX2X1_19/a_30_54# MUX2X1_19/a_2_10# INVX2_17/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1264 MUX2X1_19/a_17_10# DFFSR_1/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1265 vdd OAI21X1_0/Y MUX2X1_19/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1266 MUX2X1_19/a_30_10# OAI21X1_0/Y INVX2_17/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1267 gnd OAI21X1_0/Y MUX2X1_19/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1268 vdd DFFSR_1/D MUX2X1_19/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1269 INVX2_17/A MUX2X1_19/a_2_10# MUX2X1_19/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1270 gnd NAND2X1_2/A AOI22X1_2/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1271 INVX2_76/A DFFSR_7/S AOI22X1_2/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1272 AOI22X1_2/a_11_6# INVX2_16/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 AOI22X1_2/a_2_54# DFFSR_7/S vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1274 AOI22X1_2/a_28_6# INVX2_99/A INVX2_76/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1275 vdd INVX2_16/Y AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 INVX2_76/A INVX2_99/A AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1277 AOI22X1_2/a_2_54# NAND2X1_2/A INVX2_76/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1278 NOR2X1_37/B out_state[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1279 NAND2X1_23/a_9_6# out_state[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1280 vdd OAI21X1_21/Y NOR2X1_37/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 NOR2X1_37/B OAI21X1_21/Y NAND2X1_23/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1282 NOR2X1_9/A AOI21X1_3/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1283 NAND2X1_12/a_9_6# AOI21X1_3/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1284 vdd DFFSR_7/S NOR2X1_9/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1285 NOR2X1_9/A DFFSR_7/S NAND2X1_12/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1286 gnd OAI22X1_6/A OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1287 OAI22X1_5/a_2_6# INVX2_98/Y OAI22X1_5/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1288 OAI22X1_5/Y INVX2_80/Y OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 OAI22X1_5/Y INVX2_40/Y OAI22X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1290 OAI22X1_5/a_28_54# INVX2_80/Y OAI22X1_5/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1291 OAI22X1_5/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 OAI22X1_5/a_2_6# INVX2_40/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1293 vdd INVX2_98/Y OAI22X1_5/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1294 INVX2_14/Y INVX2_14/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1295 INVX2_14/Y INVX2_14/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1296 INVX2_25/Y INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1297 INVX2_25/Y INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1298 INVX2_69/Y INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1299 INVX2_69/Y INVX2_69/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1300 INVX2_47/Y INVX2_47/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1301 INVX2_47/Y INVX2_47/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1302 INVX2_58/Y INVX2_58/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1303 INVX2_58/Y INVX2_58/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1304 INVX2_36/Y INVX2_36/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1305 INVX2_36/Y INVX2_36/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1306 gnd INVX2_0/A XNOR2X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1307 MUX2X1_1/A INVX2_0/A XNOR2X1_8/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1308 XNOR2X1_8/a_12_41# DFFSR_7/D gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1309 XNOR2X1_8/a_18_54# XNOR2X1_8/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1310 XNOR2X1_8/a_35_6# XNOR2X1_8/a_2_6# MUX2X1_1/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1311 XNOR2X1_8/a_18_6# XNOR2X1_8/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1312 vdd INVX2_0/A XNOR2X1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1313 vdd DFFSR_7/D XNOR2X1_8/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1314 MUX2X1_1/A XNOR2X1_8/a_2_6# XNOR2X1_8/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1315 XNOR2X1_8/a_35_54# INVX2_0/A MUX2X1_1/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1316 XNOR2X1_8/a_12_41# DFFSR_7/D vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1317 gnd DFFSR_7/D XNOR2X1_8/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1318 DFFNEGX1_43/a_76_6# INVX4_0/Y DFFNEGX1_43/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1319 gnd INVX4_0/Y DFFNEGX1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1320 DFFNEGX1_43/a_66_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1321 AOI21X1_3/B DFFNEGX1_43/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1322 DFFNEGX1_43/a_23_6# INVX4_0/Y DFFNEGX1_43/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1323 DFFNEGX1_43/a_23_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1324 gnd DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1325 vdd DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1326 DFFNEGX1_43/a_61_74# DFFNEGX1_43/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1327 DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1328 DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1329 vdd AOI21X1_3/B DFFNEGX1_43/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1330 gnd AOI21X1_3/B DFFNEGX1_43/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1331 DFFNEGX1_43/a_61_6# DFFNEGX1_43/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1332 DFFNEGX1_43/a_76_84# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1333 AOI21X1_3/B DFFNEGX1_43/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1334 vdd INVX4_0/Y DFFNEGX1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1335 DFFNEGX1_43/a_31_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1336 DFFNEGX1_43/a_66_6# INVX4_0/Y DFFNEGX1_43/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1337 DFFNEGX1_43/a_17_74# INVX2_64/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1338 DFFNEGX1_43/a_31_74# INVX4_0/Y DFFNEGX1_43/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1339 DFFNEGX1_43/a_17_6# INVX2_64/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1340 DFFNEGX1_10/a_76_6# INVX2_101/Y DFFNEGX1_10/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1341 gnd INVX2_101/Y DFFNEGX1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1342 DFFNEGX1_10/a_66_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1343 INVX2_24/A DFFNEGX1_10/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1344 DFFNEGX1_10/a_23_6# INVX2_101/Y DFFNEGX1_10/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1345 DFFNEGX1_10/a_23_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1346 gnd DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1347 vdd DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1348 DFFNEGX1_10/a_61_74# DFFNEGX1_10/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1349 DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1350 DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1351 vdd INVX2_24/A DFFNEGX1_10/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1352 gnd INVX2_24/A DFFNEGX1_10/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1353 DFFNEGX1_10/a_61_6# DFFNEGX1_10/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1354 DFFNEGX1_10/a_76_84# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1355 INVX2_24/A DFFNEGX1_10/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1356 vdd INVX2_101/Y DFFNEGX1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1357 DFFNEGX1_10/a_31_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 DFFNEGX1_10/a_66_6# INVX2_101/Y DFFNEGX1_10/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1359 DFFNEGX1_10/a_17_74# OAI22X1_20/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1360 DFFNEGX1_10/a_31_74# INVX2_101/Y DFFNEGX1_10/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1361 DFFNEGX1_10/a_17_6# OAI22X1_20/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1362 DFFNEGX1_32/a_76_6# INVX4_0/Y DFFNEGX1_32/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1363 gnd INVX4_0/Y DFFNEGX1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1364 DFFNEGX1_32/a_66_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1365 INVX2_47/A DFFNEGX1_32/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1366 DFFNEGX1_32/a_23_6# INVX4_0/Y DFFNEGX1_32/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1367 DFFNEGX1_32/a_23_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1368 gnd DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1369 vdd DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1370 DFFNEGX1_32/a_61_74# DFFNEGX1_32/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1371 DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1372 DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1373 vdd INVX2_47/A DFFNEGX1_32/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1374 gnd INVX2_47/A DFFNEGX1_32/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1375 DFFNEGX1_32/a_61_6# DFFNEGX1_32/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1376 DFFNEGX1_32/a_76_84# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1377 INVX2_47/A DFFNEGX1_32/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1378 vdd INVX4_0/Y DFFNEGX1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1379 DFFNEGX1_32/a_31_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 DFFNEGX1_32/a_66_6# INVX4_0/Y DFFNEGX1_32/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1381 DFFNEGX1_32/a_17_74# OAI22X1_31/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1382 DFFNEGX1_32/a_31_74# INVX4_0/Y DFFNEGX1_32/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1383 DFFNEGX1_32/a_17_6# OAI22X1_31/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 DFFNEGX1_21/a_76_6# INVX2_102/Y DFFNEGX1_21/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1385 gnd INVX2_102/Y DFFNEGX1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1386 DFFNEGX1_21/a_66_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1387 INVX2_35/A DFFNEGX1_21/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1388 DFFNEGX1_21/a_23_6# INVX2_102/Y DFFNEGX1_21/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1389 DFFNEGX1_21/a_23_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1390 gnd DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1391 vdd DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1392 DFFNEGX1_21/a_61_74# DFFNEGX1_21/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1393 DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1394 DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1395 vdd INVX2_35/A DFFNEGX1_21/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1396 gnd INVX2_35/A DFFNEGX1_21/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1397 DFFNEGX1_21/a_61_6# DFFNEGX1_21/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1398 DFFNEGX1_21/a_76_84# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1399 INVX2_35/A DFFNEGX1_21/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1400 vdd INVX2_102/Y DFFNEGX1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1401 DFFNEGX1_21/a_31_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1402 DFFNEGX1_21/a_66_6# INVX2_102/Y DFFNEGX1_21/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1403 DFFNEGX1_21/a_17_74# OAI22X1_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1404 DFFNEGX1_21/a_31_74# INVX2_102/Y DFFNEGX1_21/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1405 DFFNEGX1_21/a_17_6# OAI22X1_10/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 gnd AOI22X1_3/C AOI22X1_3/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1407 INVX2_77/A DFFSR_7/S AOI22X1_3/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1408 AOI22X1_3/a_11_6# INVX2_17/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 AOI22X1_3/a_2_54# DFFSR_7/S vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1410 AOI22X1_3/a_28_6# INVX2_99/A INVX2_77/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1411 vdd INVX2_17/Y AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1412 INVX2_77/A INVX2_99/A AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1413 AOI22X1_3/a_2_54# AOI22X1_3/C INVX2_77/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1414 OAI21X1_21/C in_enter vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1415 NAND2X1_24/a_9_6# in_enter gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1416 vdd INVX2_63/Y OAI21X1_21/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1417 OAI21X1_21/C INVX2_63/Y NAND2X1_24/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1418 XNOR2X1_22/A XOR2X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1419 NAND2X1_13/a_9_6# XOR2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1420 vdd XOR2X1_3/B XNOR2X1_22/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1421 XNOR2X1_22/A XOR2X1_3/B NAND2X1_13/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1422 gnd OAI22X1_6/A OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1423 OAI22X1_6/a_2_6# INVX2_98/Y OAI22X1_6/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1424 OAI22X1_6/Y INVX2_81/Y OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1425 OAI22X1_6/Y INVX2_39/Y OAI22X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1426 OAI22X1_6/a_28_54# INVX2_81/Y OAI22X1_6/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1427 OAI22X1_6/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 OAI22X1_6/a_2_6# INVX2_39/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 vdd INVX2_98/Y OAI22X1_6/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 INVX2_15/Y INVX2_15/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1431 INVX2_15/Y INVX2_15/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1432 INVX2_26/Y INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1433 INVX2_26/Y INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1434 INVX2_37/Y INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1435 INVX2_37/Y INVX2_37/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1436 out_Bnum[2] INVX2_59/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1437 out_Bnum[2] INVX2_59/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1438 INVX2_48/Y INVX2_48/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1439 INVX2_48/Y INVX2_48/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1440 gnd INVX2_1/A XNOR2X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1441 MUX2X1_0/A INVX2_1/A XNOR2X1_9/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1442 XNOR2X1_9/a_12_41# NOR2X1_5/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1443 XNOR2X1_9/a_18_54# XNOR2X1_9/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1444 XNOR2X1_9/a_35_6# XNOR2X1_9/a_2_6# MUX2X1_0/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1445 XNOR2X1_9/a_18_6# XNOR2X1_9/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 vdd INVX2_1/A XNOR2X1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1447 vdd NOR2X1_5/A XNOR2X1_9/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1448 MUX2X1_0/A XNOR2X1_9/a_2_6# XNOR2X1_9/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1449 XNOR2X1_9/a_35_54# INVX2_1/A MUX2X1_0/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1450 XNOR2X1_9/a_12_41# NOR2X1_5/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1451 gnd NOR2X1_5/A XNOR2X1_9/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 DFFNEGX1_44/a_76_6# INVX4_0/Y DFFNEGX1_44/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1453 gnd INVX4_0/Y DFFNEGX1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1454 DFFNEGX1_44/a_66_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1455 INVX2_99/A DFFNEGX1_44/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1456 DFFNEGX1_44/a_23_6# INVX4_0/Y DFFNEGX1_44/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1457 DFFNEGX1_44/a_23_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1458 gnd DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1459 vdd DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1460 DFFNEGX1_44/a_61_74# DFFNEGX1_44/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1461 DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1462 DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1463 vdd INVX2_99/A DFFNEGX1_44/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1464 gnd INVX2_99/A DFFNEGX1_44/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1465 DFFNEGX1_44/a_61_6# DFFNEGX1_44/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1466 DFFNEGX1_44/a_76_84# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1467 INVX2_99/A DFFNEGX1_44/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1468 vdd INVX4_0/Y DFFNEGX1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1469 DFFNEGX1_44/a_31_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1470 DFFNEGX1_44/a_66_6# INVX4_0/Y DFFNEGX1_44/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1471 DFFNEGX1_44/a_17_74# INVX2_62/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 DFFNEGX1_44/a_31_74# INVX4_0/Y DFFNEGX1_44/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 DFFNEGX1_44/a_17_6# INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1474 DFFNEGX1_11/a_76_6# INVX2_101/Y DFFNEGX1_11/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1475 gnd INVX2_101/Y DFFNEGX1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1476 DFFNEGX1_11/a_66_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1477 INVX2_25/A DFFNEGX1_11/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1478 DFFNEGX1_11/a_23_6# INVX2_101/Y DFFNEGX1_11/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1479 DFFNEGX1_11/a_23_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1480 gnd DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1481 vdd DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1482 DFFNEGX1_11/a_61_74# DFFNEGX1_11/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1483 DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1484 DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1485 vdd INVX2_25/A DFFNEGX1_11/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1486 gnd INVX2_25/A DFFNEGX1_11/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1487 DFFNEGX1_11/a_61_6# DFFNEGX1_11/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1488 DFFNEGX1_11/a_76_84# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1489 INVX2_25/A DFFNEGX1_11/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1490 vdd INVX2_101/Y DFFNEGX1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1491 DFFNEGX1_11/a_31_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1492 DFFNEGX1_11/a_66_6# INVX2_101/Y DFFNEGX1_11/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1493 DFFNEGX1_11/a_17_74# OAI22X1_19/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 DFFNEGX1_11/a_31_74# INVX2_101/Y DFFNEGX1_11/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1495 DFFNEGX1_11/a_17_6# OAI22X1_19/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 DFFNEGX1_33/a_76_6# INVX4_0/Y DFFNEGX1_33/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1497 gnd INVX4_0/Y DFFNEGX1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1498 DFFNEGX1_33/a_66_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1499 INVX2_49/A DFFNEGX1_33/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1500 DFFNEGX1_33/a_23_6# INVX4_0/Y DFFNEGX1_33/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1501 DFFNEGX1_33/a_23_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1502 gnd DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1503 vdd DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1504 DFFNEGX1_33/a_61_74# DFFNEGX1_33/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1505 DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1506 DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1507 vdd INVX2_49/A DFFNEGX1_33/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1508 gnd INVX2_49/A DFFNEGX1_33/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1509 DFFNEGX1_33/a_61_6# DFFNEGX1_33/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1510 DFFNEGX1_33/a_76_84# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1511 INVX2_49/A DFFNEGX1_33/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1512 vdd INVX4_0/Y DFFNEGX1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1513 DFFNEGX1_33/a_31_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1514 DFFNEGX1_33/a_66_6# INVX4_0/Y DFFNEGX1_33/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1515 DFFNEGX1_33/a_17_74# OAI22X1_30/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1516 DFFNEGX1_33/a_31_74# INVX4_0/Y DFFNEGX1_33/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 DFFNEGX1_33/a_17_6# OAI22X1_30/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 DFFNEGX1_22/a_76_6# INVX2_102/Y DFFNEGX1_22/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1519 gnd INVX2_102/Y DFFNEGX1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1520 DFFNEGX1_22/a_66_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1521 INVX2_36/A DFFNEGX1_22/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1522 DFFNEGX1_22/a_23_6# INVX2_102/Y DFFNEGX1_22/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1523 DFFNEGX1_22/a_23_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1524 gnd DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1525 vdd DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1526 DFFNEGX1_22/a_61_74# DFFNEGX1_22/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1527 DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1528 DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1529 vdd INVX2_36/A DFFNEGX1_22/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1530 gnd INVX2_36/A DFFNEGX1_22/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1531 DFFNEGX1_22/a_61_6# DFFNEGX1_22/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1532 DFFNEGX1_22/a_76_84# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1533 INVX2_36/A DFFNEGX1_22/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1534 vdd INVX2_102/Y DFFNEGX1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1535 DFFNEGX1_22/a_31_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 DFFNEGX1_22/a_66_6# INVX2_102/Y DFFNEGX1_22/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1537 DFFNEGX1_22/a_17_74# OAI22X1_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1538 DFFNEGX1_22/a_31_74# INVX2_102/Y DFFNEGX1_22/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1539 DFFNEGX1_22/a_17_6# OAI22X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1540 gnd XOR2X1_4/A AOI22X1_4/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1541 INVX2_58/A XOR2X1_5/B AOI22X1_4/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1542 AOI22X1_4/a_11_6# XOR2X1_5/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1543 AOI22X1_4/a_2_54# XOR2X1_5/B vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1544 AOI22X1_4/a_28_6# XOR2X1_5/Y INVX2_58/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1545 vdd XOR2X1_5/A AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1546 INVX2_58/A XOR2X1_5/Y AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1547 AOI22X1_4/a_2_54# XOR2X1_4/A INVX2_58/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1548 OAI21X1_17/B XNOR2X1_32/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1549 NAND2X1_14/a_9_6# XNOR2X1_32/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1550 vdd XNOR2X1_31/Y OAI21X1_17/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1551 OAI21X1_17/B XNOR2X1_31/Y NAND2X1_14/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1552 gnd INVX2_67/A OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1553 OAI22X1_7/a_2_6# INVX2_67/Y OAI22X1_7/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1554 OAI22X1_7/Y OAI22X1_7/D OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1555 OAI22X1_7/Y INVX2_38/Y OAI22X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1556 OAI22X1_7/a_28_54# OAI22X1_7/D OAI22X1_7/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1557 OAI22X1_7/a_9_54# INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 OAI22X1_7/a_2_6# INVX2_38/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1559 vdd INVX2_67/Y OAI22X1_7/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1560 INVX2_16/Y INVX2_16/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1561 INVX2_16/Y INVX2_16/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1562 INVX2_27/Y INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1563 INVX2_27/Y INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1564 INVX2_38/Y INVX2_38/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1565 INVX2_38/Y INVX2_38/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1566 INVX2_49/Y INVX2_49/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1567 INVX2_49/Y INVX2_49/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1568 gnd MUX2X1_0/A MUX2X1_0/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1569 MUX2X1_0/a_17_50# INVX2_1/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1570 MUX2X1_0/Y NOR2X1_5/Y MUX2X1_0/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1571 MUX2X1_0/a_30_54# MUX2X1_0/a_2_10# MUX2X1_0/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1572 MUX2X1_0/a_17_10# INVX2_1/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1573 vdd NOR2X1_5/Y MUX2X1_0/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1574 MUX2X1_0/a_30_10# NOR2X1_5/Y MUX2X1_0/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1575 gnd NOR2X1_5/Y MUX2X1_0/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1576 vdd MUX2X1_0/A MUX2X1_0/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 MUX2X1_0/Y MUX2X1_0/a_2_10# MUX2X1_0/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 DFFNEGX1_23/a_76_6# INVX2_102/Y DFFNEGX1_23/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1579 gnd INVX2_102/Y DFFNEGX1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1580 DFFNEGX1_23/a_66_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1581 INVX2_37/A DFFNEGX1_23/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1582 DFFNEGX1_23/a_23_6# INVX2_102/Y DFFNEGX1_23/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1583 DFFNEGX1_23/a_23_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1584 gnd DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1585 vdd DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1586 DFFNEGX1_23/a_61_74# DFFNEGX1_23/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1587 DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1588 DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1589 vdd INVX2_37/A DFFNEGX1_23/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1590 gnd INVX2_37/A DFFNEGX1_23/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1591 DFFNEGX1_23/a_61_6# DFFNEGX1_23/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1592 DFFNEGX1_23/a_76_84# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1593 INVX2_37/A DFFNEGX1_23/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1594 vdd INVX2_102/Y DFFNEGX1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1595 DFFNEGX1_23/a_31_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 DFFNEGX1_23/a_66_6# INVX2_102/Y DFFNEGX1_23/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1597 DFFNEGX1_23/a_17_74# OAI22X1_8/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1598 DFFNEGX1_23/a_31_74# INVX2_102/Y DFFNEGX1_23/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1599 DFFNEGX1_23/a_17_6# OAI22X1_8/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1600 DFFNEGX1_12/a_76_6# INVX2_101/Y DFFNEGX1_12/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1601 gnd INVX2_101/Y DFFNEGX1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1602 DFFNEGX1_12/a_66_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1603 INVX2_26/A DFFNEGX1_12/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1604 DFFNEGX1_12/a_23_6# INVX2_101/Y DFFNEGX1_12/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1605 DFFNEGX1_12/a_23_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1606 gnd DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1607 vdd DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1608 DFFNEGX1_12/a_61_74# DFFNEGX1_12/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1609 DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1610 DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1611 vdd INVX2_26/A DFFNEGX1_12/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1612 gnd INVX2_26/A DFFNEGX1_12/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 DFFNEGX1_12/a_61_6# DFFNEGX1_12/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1614 DFFNEGX1_12/a_76_84# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1615 INVX2_26/A DFFNEGX1_12/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1616 vdd INVX2_101/Y DFFNEGX1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1617 DFFNEGX1_12/a_31_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1618 DFFNEGX1_12/a_66_6# INVX2_101/Y DFFNEGX1_12/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1619 DFFNEGX1_12/a_17_74# OAI22X1_18/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1620 DFFNEGX1_12/a_31_74# INVX2_101/Y DFFNEGX1_12/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 DFFNEGX1_12/a_17_6# OAI22X1_18/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1622 DFFNEGX1_34/a_76_6# INVX4_0/Y DFFNEGX1_34/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1623 gnd INVX4_0/Y DFFNEGX1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1624 DFFNEGX1_34/a_66_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1625 INVX2_50/A DFFNEGX1_34/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1626 DFFNEGX1_34/a_23_6# INVX4_0/Y DFFNEGX1_34/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1627 DFFNEGX1_34/a_23_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1628 gnd DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1629 vdd DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1630 DFFNEGX1_34/a_61_74# DFFNEGX1_34/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1631 DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1632 DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1633 vdd INVX2_50/A DFFNEGX1_34/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1634 gnd INVX2_50/A DFFNEGX1_34/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1635 DFFNEGX1_34/a_61_6# DFFNEGX1_34/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1636 DFFNEGX1_34/a_76_84# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1637 INVX2_50/A DFFNEGX1_34/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1638 vdd INVX4_0/Y DFFNEGX1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1639 DFFNEGX1_34/a_31_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1640 DFFNEGX1_34/a_66_6# INVX4_0/Y DFFNEGX1_34/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1641 DFFNEGX1_34/a_17_74# OAI22X1_29/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1642 DFFNEGX1_34/a_31_74# INVX4_0/Y DFFNEGX1_34/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1643 DFFNEGX1_34/a_17_6# OAI22X1_29/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1644 OAI21X1_8/C INVX2_73/Y vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1645 NAND3X1_0/a_9_6# INVX2_73/Y gnd Gnd nfet w=30 l=2
+  ad=45p pd=33u as=0.15n ps=70u
M1646 OAI21X1_8/C NOR2X1_7/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1647 OAI21X1_8/C NOR2X1_7/Y NAND3X1_0/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=45p ps=33u
M1648 vdd NOR2X1_9/Y OAI21X1_8/C vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1649 NAND3X1_0/a_14_6# NOR2X1_9/Y NAND3X1_0/a_9_6# Gnd nfet w=30 l=2
+  ad=45p pd=33u as=45p ps=33u
M1650 gnd NOR2X1_16/Y AOI22X1_5/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1651 AOI22X1_5/Y NOR2X1_17/Y AOI22X1_5/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1652 AOI22X1_5/a_11_6# NOR2X1_18/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1653 AOI22X1_5/a_2_54# NOR2X1_17/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1654 AOI22X1_5/a_28_6# NOR2X1_15/Y AOI22X1_5/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1655 vdd NOR2X1_18/Y AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1656 AOI22X1_5/Y NOR2X1_15/Y AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1657 AOI22X1_5/a_2_54# NOR2X1_16/Y AOI22X1_5/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1658 OAI21X1_17/A XNOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1659 NAND2X1_15/a_9_6# XNOR2X1_34/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1660 vdd XNOR2X1_33/Y OAI21X1_17/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 OAI21X1_17/A XNOR2X1_33/Y NAND2X1_15/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1662 gnd INVX2_37/A XNOR2X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1663 XNOR2X1_90/Y INVX2_37/A XNOR2X1_90/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1664 XNOR2X1_90/a_12_41# INVX2_41/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1665 XNOR2X1_90/a_18_54# XNOR2X1_90/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1666 XNOR2X1_90/a_35_6# XNOR2X1_90/a_2_6# XNOR2X1_90/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1667 XNOR2X1_90/a_18_6# XNOR2X1_90/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1668 vdd INVX2_37/A XNOR2X1_90/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1669 vdd INVX2_41/A XNOR2X1_90/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1670 XNOR2X1_90/Y XNOR2X1_90/a_2_6# XNOR2X1_90/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1671 XNOR2X1_90/a_35_54# INVX2_37/A XNOR2X1_90/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1672 XNOR2X1_90/a_12_41# INVX2_41/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1673 gnd INVX2_41/A XNOR2X1_90/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1674 gnd INVX2_67/A OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1675 OAI22X1_8/a_2_6# INVX2_67/Y OAI22X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1676 OAI22X1_8/Y OAI22X1_8/D OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 OAI22X1_8/Y INVX2_37/Y OAI22X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1678 OAI22X1_8/a_28_54# OAI22X1_8/D OAI22X1_8/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1679 OAI22X1_8/a_9_54# INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 OAI22X1_8/a_2_6# INVX2_37/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1681 vdd INVX2_67/Y OAI22X1_8/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1682 INVX2_17/Y INVX2_17/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1683 INVX2_17/Y INVX2_17/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1684 INVX2_28/Y INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1685 INVX2_28/Y INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1686 INVX2_39/Y INVX2_39/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1687 INVX2_39/Y INVX2_39/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1688 gnd XOR2X1_2/Y XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=100p ps=50u
M1689 DFFSR_0/D XOR2X1_0/a_2_6# XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M1690 XOR2X1_0/a_13_43# XOR2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=70p ps=27u
M1691 XOR2X1_0/a_18_54# XOR2X1_0/a_13_43# vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.14n ps=47u
M1692 XOR2X1_0/a_35_6# XOR2X1_2/Y DFFSR_0/D Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M1693 XOR2X1_0/a_18_6# XOR2X1_0/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=70p ps=27u
M1694 vdd XOR2X1_2/Y XOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=0.2n ps=90u
M1695 vdd XOR2X1_1/Y XOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=59.999996p ps=43u
M1696 DFFSR_0/D XOR2X1_2/Y XOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=0.2n pd=50u as=59.999996p ps=43u
M1697 XOR2X1_0/a_35_54# XOR2X1_0/a_2_6# DFFSR_0/D vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=50u
M1698 XOR2X1_0/a_13_43# XOR2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.14n ps=47u
M1699 gnd XOR2X1_1/Y XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=29.999998p ps=23u
M1700 gnd MUX2X1_1/A MUX2X1_1/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1701 MUX2X1_1/a_17_50# DFFSR_7/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1702 INVX2_2/A NOR2X1_5/Y MUX2X1_1/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1703 MUX2X1_1/a_30_54# MUX2X1_1/a_2_10# INVX2_2/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1704 MUX2X1_1/a_17_10# DFFSR_7/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1705 vdd NOR2X1_5/Y MUX2X1_1/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1706 MUX2X1_1/a_30_10# NOR2X1_5/Y INVX2_2/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1707 gnd NOR2X1_5/Y MUX2X1_1/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1708 vdd MUX2X1_1/A MUX2X1_1/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1709 INVX2_2/A MUX2X1_1/a_2_10# MUX2X1_1/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1710 DFFNEGX1_13/a_76_6# INVX2_102/Y DFFNEGX1_13/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1711 gnd INVX2_102/Y DFFNEGX1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1712 DFFNEGX1_13/a_66_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1713 INVX2_27/A DFFNEGX1_13/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1714 DFFNEGX1_13/a_23_6# INVX2_102/Y DFFNEGX1_13/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1715 DFFNEGX1_13/a_23_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1716 gnd DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1717 vdd DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1718 DFFNEGX1_13/a_61_74# DFFNEGX1_13/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1719 DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1720 DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1721 vdd INVX2_27/A DFFNEGX1_13/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1722 gnd INVX2_27/A DFFNEGX1_13/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1723 DFFNEGX1_13/a_61_6# DFFNEGX1_13/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1724 DFFNEGX1_13/a_76_84# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1725 INVX2_27/A DFFNEGX1_13/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1726 vdd INVX2_102/Y DFFNEGX1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1727 DFFNEGX1_13/a_31_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1728 DFFNEGX1_13/a_66_6# INVX2_102/Y DFFNEGX1_13/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1729 DFFNEGX1_13/a_17_74# OAI22X1_14/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1730 DFFNEGX1_13/a_31_74# INVX2_102/Y DFFNEGX1_13/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1731 DFFNEGX1_13/a_17_6# OAI22X1_14/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1732 DFFNEGX1_24/a_76_6# INVX2_102/Y DFFNEGX1_24/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1733 gnd INVX2_102/Y DFFNEGX1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1734 DFFNEGX1_24/a_66_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1735 INVX2_38/A DFFNEGX1_24/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1736 DFFNEGX1_24/a_23_6# INVX2_102/Y DFFNEGX1_24/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1737 DFFNEGX1_24/a_23_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1738 gnd DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1739 vdd DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1740 DFFNEGX1_24/a_61_74# DFFNEGX1_24/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1741 DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1742 DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1743 vdd INVX2_38/A DFFNEGX1_24/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1744 gnd INVX2_38/A DFFNEGX1_24/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1745 DFFNEGX1_24/a_61_6# DFFNEGX1_24/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1746 DFFNEGX1_24/a_76_84# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1747 INVX2_38/A DFFNEGX1_24/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1748 vdd INVX2_102/Y DFFNEGX1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1749 DFFNEGX1_24/a_31_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1750 DFFNEGX1_24/a_66_6# INVX2_102/Y DFFNEGX1_24/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1751 DFFNEGX1_24/a_17_74# OAI22X1_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1752 DFFNEGX1_24/a_31_74# INVX2_102/Y DFFNEGX1_24/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1753 DFFNEGX1_24/a_17_6# OAI22X1_7/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1754 DFFNEGX1_35/a_76_6# INVX4_0/Y DFFNEGX1_35/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1755 gnd INVX4_0/Y DFFNEGX1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1756 DFFNEGX1_35/a_66_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1757 INVX2_51/A DFFNEGX1_35/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1758 DFFNEGX1_35/a_23_6# INVX4_0/Y DFFNEGX1_35/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1759 DFFNEGX1_35/a_23_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1760 gnd DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1761 vdd DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1762 DFFNEGX1_35/a_61_74# DFFNEGX1_35/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1763 DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1764 DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1765 vdd INVX2_51/A DFFNEGX1_35/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1766 gnd INVX2_51/A DFFNEGX1_35/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1767 DFFNEGX1_35/a_61_6# DFFNEGX1_35/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1768 DFFNEGX1_35/a_76_84# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1769 INVX2_51/A DFFNEGX1_35/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1770 vdd INVX4_0/Y DFFNEGX1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1771 DFFNEGX1_35/a_31_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1772 DFFNEGX1_35/a_66_6# INVX4_0/Y DFFNEGX1_35/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1773 DFFNEGX1_35/a_17_74# OAI22X1_28/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1774 DFFNEGX1_35/a_31_74# INVX4_0/Y DFFNEGX1_35/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1775 DFFNEGX1_35/a_17_6# OAI22X1_28/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1776 OAI21X1_9/C INVX2_72/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M1777 NAND3X1_1/a_9_6# INVX2_72/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M1778 OAI21X1_9/C INVX2_73/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1779 OAI21X1_9/C INVX2_73/Y NAND3X1_1/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M1780 vdd NOR2X1_7/A OAI21X1_9/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1781 NAND3X1_1/a_14_6# NOR2X1_7/A NAND3X1_1/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1782 gnd NOR2X1_20/Y AOI22X1_6/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1783 AOI22X1_6/Y NOR2X1_21/Y AOI22X1_6/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1784 AOI22X1_6/a_11_6# NOR2X1_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1785 AOI22X1_6/a_2_54# NOR2X1_21/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1786 AOI22X1_6/a_28_6# NOR2X1_19/Y AOI22X1_6/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1787 vdd NOR2X1_22/Y AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1788 AOI22X1_6/Y NOR2X1_19/Y AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1789 AOI22X1_6/a_2_54# NOR2X1_20/Y AOI22X1_6/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1790 OAI21X1_18/B XNOR2X1_44/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1791 NAND2X1_16/a_9_6# XNOR2X1_44/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1792 vdd XNOR2X1_43/Y OAI21X1_18/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1793 OAI21X1_18/B XNOR2X1_43/Y NAND2X1_16/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1794 gnd INVX2_54/Y XNOR2X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1795 NOR2X1_32/A INVX2_54/Y XNOR2X1_80/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1796 XNOR2X1_80/a_12_41# INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1797 XNOR2X1_80/a_18_54# XNOR2X1_80/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1798 XNOR2X1_80/a_35_6# XNOR2X1_80/a_2_6# NOR2X1_32/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1799 XNOR2X1_80/a_18_6# XNOR2X1_80/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1800 vdd INVX2_54/Y XNOR2X1_80/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1801 vdd INVX2_30/A XNOR2X1_80/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1802 NOR2X1_32/A XNOR2X1_80/a_2_6# XNOR2X1_80/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1803 XNOR2X1_80/a_35_54# INVX2_54/Y NOR2X1_32/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1804 XNOR2X1_80/a_12_41# INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1805 gnd INVX2_30/A XNOR2X1_80/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1806 gnd INVX2_67/A OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1807 OAI22X1_9/a_2_6# INVX2_67/Y OAI22X1_9/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1808 OAI22X1_9/Y OAI22X1_9/D OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1809 OAI22X1_9/Y INVX2_36/Y OAI22X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1810 OAI22X1_9/a_28_54# OAI22X1_9/D OAI22X1_9/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1811 OAI22X1_9/a_9_54# INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1812 OAI22X1_9/a_2_6# INVX2_36/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1813 vdd INVX2_67/Y OAI22X1_9/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1814 INVX2_29/Y INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1815 INVX2_29/Y INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1816 INVX2_18/Y INVX2_18/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1817 INVX2_18/Y INVX2_18/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1818 gnd DFFSR_5/D XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1819 XOR2X1_1/Y XOR2X1_1/a_2_6# XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1820 XOR2X1_1/a_13_43# DFFSR_4/D gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1821 XOR2X1_1/a_18_54# XOR2X1_1/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1822 XOR2X1_1/a_35_6# DFFSR_5/D XOR2X1_1/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1823 XOR2X1_1/a_18_6# XOR2X1_1/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1824 vdd DFFSR_5/D XOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1825 vdd DFFSR_4/D XOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1826 XOR2X1_1/Y DFFSR_5/D XOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1827 XOR2X1_1/a_35_54# XOR2X1_1/a_2_6# XOR2X1_1/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1828 XOR2X1_1/a_13_43# DFFSR_4/D vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1829 gnd DFFSR_4/D XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1830 gnd INVX2_0/Y MUX2X1_2/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1831 MUX2X1_2/a_17_50# INVX2_0/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1832 INVX2_3/A NOR2X1_5/Y MUX2X1_2/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1833 MUX2X1_2/a_30_54# MUX2X1_2/a_2_10# INVX2_3/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1834 MUX2X1_2/a_17_10# INVX2_0/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1835 vdd NOR2X1_5/Y MUX2X1_2/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1836 MUX2X1_2/a_30_10# NOR2X1_5/Y INVX2_3/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1837 gnd NOR2X1_5/Y MUX2X1_2/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1838 vdd INVX2_0/Y MUX2X1_2/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1839 INVX2_3/A MUX2X1_2/a_2_10# MUX2X1_2/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1840 DFFNEGX1_14/a_76_6# INVX2_102/Y DFFNEGX1_14/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1841 gnd INVX2_102/Y DFFNEGX1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1842 DFFNEGX1_14/a_66_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1843 INVX2_28/A DFFNEGX1_14/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1844 DFFNEGX1_14/a_23_6# INVX2_102/Y DFFNEGX1_14/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1845 DFFNEGX1_14/a_23_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1846 gnd DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1847 vdd DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1848 DFFNEGX1_14/a_61_74# DFFNEGX1_14/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1849 DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1850 DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1851 vdd INVX2_28/A DFFNEGX1_14/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1852 gnd INVX2_28/A DFFNEGX1_14/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1853 DFFNEGX1_14/a_61_6# DFFNEGX1_14/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1854 DFFNEGX1_14/a_76_84# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1855 INVX2_28/A DFFNEGX1_14/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1856 vdd INVX2_102/Y DFFNEGX1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1857 DFFNEGX1_14/a_31_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1858 DFFNEGX1_14/a_66_6# INVX2_102/Y DFFNEGX1_14/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1859 DFFNEGX1_14/a_17_74# OAI22X1_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1860 DFFNEGX1_14/a_31_74# INVX2_102/Y DFFNEGX1_14/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1861 DFFNEGX1_14/a_17_6# OAI22X1_13/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1862 DFFNEGX1_36/a_76_6# INVX4_0/Y DFFNEGX1_36/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1863 gnd INVX4_0/Y DFFNEGX1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1864 DFFNEGX1_36/a_66_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1865 INVX2_52/A DFFNEGX1_36/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1866 DFFNEGX1_36/a_23_6# INVX4_0/Y DFFNEGX1_36/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1867 DFFNEGX1_36/a_23_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1868 gnd DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1869 vdd DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1870 DFFNEGX1_36/a_61_74# DFFNEGX1_36/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1871 DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1872 DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1873 vdd INVX2_52/A DFFNEGX1_36/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1874 gnd INVX2_52/A DFFNEGX1_36/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1875 DFFNEGX1_36/a_61_6# DFFNEGX1_36/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1876 DFFNEGX1_36/a_76_84# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1877 INVX2_52/A DFFNEGX1_36/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1878 vdd INVX4_0/Y DFFNEGX1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1879 DFFNEGX1_36/a_31_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1880 DFFNEGX1_36/a_66_6# INVX4_0/Y DFFNEGX1_36/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1881 DFFNEGX1_36/a_17_74# OAI22X1_27/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1882 DFFNEGX1_36/a_31_74# INVX4_0/Y DFFNEGX1_36/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1883 DFFNEGX1_36/a_17_6# OAI22X1_27/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1884 DFFNEGX1_25/a_76_6# INVX4_0/Y DFFNEGX1_25/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1885 gnd INVX4_0/Y DFFNEGX1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1886 DFFNEGX1_25/a_66_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1887 INVX2_39/A DFFNEGX1_25/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1888 DFFNEGX1_25/a_23_6# INVX4_0/Y DFFNEGX1_25/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1889 DFFNEGX1_25/a_23_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1890 gnd DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1891 vdd DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1892 DFFNEGX1_25/a_61_74# DFFNEGX1_25/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1893 DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1894 DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1895 vdd INVX2_39/A DFFNEGX1_25/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1896 gnd INVX2_39/A DFFNEGX1_25/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1897 DFFNEGX1_25/a_61_6# DFFNEGX1_25/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1898 DFFNEGX1_25/a_76_84# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1899 INVX2_39/A DFFNEGX1_25/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1900 vdd INVX4_0/Y DFFNEGX1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1901 DFFNEGX1_25/a_31_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1902 DFFNEGX1_25/a_66_6# INVX4_0/Y DFFNEGX1_25/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1903 DFFNEGX1_25/a_17_74# OAI22X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1904 DFFNEGX1_25/a_31_74# INVX4_0/Y DFFNEGX1_25/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1905 DFFNEGX1_25/a_17_6# OAI22X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1906 NAND3X1_2/Y INVX2_72/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M1907 NAND3X1_2/a_9_6# INVX2_72/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M1908 NAND3X1_2/Y INVX2_73/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1909 NAND3X1_2/Y INVX2_73/Y NAND3X1_2/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M1910 vdd NOR2X1_14/Y NAND3X1_2/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1911 NAND3X1_2/a_14_6# NOR2X1_14/Y NAND3X1_2/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M1912 gnd NOR2X1_24/Y AOI22X1_7/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1913 AOI22X1_7/Y NOR2X1_25/Y AOI22X1_7/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1914 AOI22X1_7/a_11_6# NOR2X1_26/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1915 AOI22X1_7/a_2_54# NOR2X1_25/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1916 AOI22X1_7/a_28_6# NOR2X1_23/Y AOI22X1_7/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1917 vdd NOR2X1_26/Y AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1918 AOI22X1_7/Y NOR2X1_23/Y AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1919 AOI22X1_7/a_2_54# NOR2X1_24/Y AOI22X1_7/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1920 OAI21X1_18/A XNOR2X1_46/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1921 NAND2X1_17/a_9_6# XNOR2X1_46/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1922 vdd XNOR2X1_45/Y OAI21X1_18/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1923 OAI21X1_18/A XNOR2X1_45/Y NAND2X1_17/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1924 gnd INVX2_52/A XNOR2X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1925 XNOR2X1_70/Y INVX2_52/A XNOR2X1_70/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1926 XNOR2X1_70/a_12_41# INVX2_23/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1927 XNOR2X1_70/a_18_54# XNOR2X1_70/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1928 XNOR2X1_70/a_35_6# XNOR2X1_70/a_2_6# XNOR2X1_70/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1929 XNOR2X1_70/a_18_6# XNOR2X1_70/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1930 vdd INVX2_52/A XNOR2X1_70/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1931 vdd INVX2_23/A XNOR2X1_70/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1932 XNOR2X1_70/Y XNOR2X1_70/a_2_6# XNOR2X1_70/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1933 XNOR2X1_70/a_35_54# INVX2_52/A XNOR2X1_70/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1934 XNOR2X1_70/a_12_41# INVX2_23/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1935 gnd INVX2_23/A XNOR2X1_70/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1936 gnd INVX2_55/A XNOR2X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1937 XNOR2X1_81/Y INVX2_55/A XNOR2X1_81/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1938 XNOR2X1_81/a_12_41# INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1939 XNOR2X1_81/a_18_54# XNOR2X1_81/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1940 XNOR2X1_81/a_35_6# XNOR2X1_81/a_2_6# XNOR2X1_81/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1941 XNOR2X1_81/a_18_6# XNOR2X1_81/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1942 vdd INVX2_55/A XNOR2X1_81/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1943 vdd INVX2_29/A XNOR2X1_81/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1944 XNOR2X1_81/Y XNOR2X1_81/a_2_6# XNOR2X1_81/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1945 XNOR2X1_81/a_35_54# INVX2_55/A XNOR2X1_81/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1946 XNOR2X1_81/a_12_41# INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1947 gnd INVX2_29/A XNOR2X1_81/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1948 NOR2X1_7/A INVX2_19/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1949 NOR2X1_7/A INVX2_19/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1950 gnd INVX2_1/A XOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1951 XOR2X1_2/Y XOR2X1_2/a_2_6# XOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1952 XOR2X1_2/a_13_43# INVX2_0/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1953 XOR2X1_2/a_18_54# XOR2X1_2/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1954 XOR2X1_2/a_35_6# INVX2_1/A XOR2X1_2/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1955 XOR2X1_2/a_18_6# XOR2X1_2/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1956 vdd INVX2_1/A XOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1957 vdd INVX2_0/A XOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1958 XOR2X1_2/Y INVX2_1/A XOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1959 XOR2X1_2/a_35_54# XOR2X1_2/a_2_6# XOR2X1_2/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 XOR2X1_2/a_13_43# INVX2_0/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1961 gnd INVX2_0/A XOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1962 gnd DFFSR_5/D MUX2X1_3/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1963 MUX2X1_3/a_17_50# DFFSR_5/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1964 INVX2_4/A NOR2X1_5/Y MUX2X1_3/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1965 MUX2X1_3/a_30_54# MUX2X1_3/a_2_10# INVX2_4/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1966 MUX2X1_3/a_17_10# DFFSR_5/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1967 vdd NOR2X1_5/Y MUX2X1_3/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1968 MUX2X1_3/a_30_10# NOR2X1_5/Y INVX2_4/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1969 gnd NOR2X1_5/Y MUX2X1_3/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1970 vdd DFFSR_5/D MUX2X1_3/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1971 INVX2_4/A MUX2X1_3/a_2_10# MUX2X1_3/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1972 DFFNEGX1_15/a_76_6# INVX2_102/Y DFFNEGX1_15/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1973 gnd INVX2_102/Y DFFNEGX1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1974 DFFNEGX1_15/a_66_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1975 INVX2_29/A DFFNEGX1_15/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1976 DFFNEGX1_15/a_23_6# INVX2_102/Y DFFNEGX1_15/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1977 DFFNEGX1_15/a_23_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1978 gnd DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1979 vdd DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1980 DFFNEGX1_15/a_61_74# DFFNEGX1_15/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1981 DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1982 DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1983 vdd INVX2_29/A DFFNEGX1_15/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1984 gnd INVX2_29/A DFFNEGX1_15/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1985 DFFNEGX1_15/a_61_6# DFFNEGX1_15/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1986 DFFNEGX1_15/a_76_84# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1987 INVX2_29/A DFFNEGX1_15/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1988 vdd INVX2_102/Y DFFNEGX1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1989 DFFNEGX1_15/a_31_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1990 DFFNEGX1_15/a_66_6# INVX2_102/Y DFFNEGX1_15/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1991 DFFNEGX1_15/a_17_74# OAI22X1_12/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1992 DFFNEGX1_15/a_31_74# INVX2_102/Y DFFNEGX1_15/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1993 DFFNEGX1_15/a_17_6# OAI22X1_12/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1994 DFFNEGX1_37/a_76_6# INVX4_0/Y DFFNEGX1_37/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1995 gnd INVX4_0/Y DFFNEGX1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1996 DFFNEGX1_37/a_66_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1997 INVX2_54/A DFFNEGX1_37/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1998 DFFNEGX1_37/a_23_6# INVX4_0/Y DFFNEGX1_37/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1999 DFFNEGX1_37/a_23_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2000 gnd DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2001 vdd DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2002 DFFNEGX1_37/a_61_74# DFFNEGX1_37/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2003 DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2004 DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2005 vdd INVX2_54/A DFFNEGX1_37/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2006 gnd INVX2_54/A DFFNEGX1_37/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2007 DFFNEGX1_37/a_61_6# DFFNEGX1_37/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2008 DFFNEGX1_37/a_76_84# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2009 INVX2_54/A DFFNEGX1_37/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2010 vdd INVX4_0/Y DFFNEGX1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2011 DFFNEGX1_37/a_31_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2012 DFFNEGX1_37/a_66_6# INVX4_0/Y DFFNEGX1_37/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2013 DFFNEGX1_37/a_17_74# OAI22X1_26/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2014 DFFNEGX1_37/a_31_74# INVX4_0/Y DFFNEGX1_37/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2015 DFFNEGX1_37/a_17_6# OAI22X1_26/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2016 DFFNEGX1_26/a_76_6# INVX4_0/Y DFFNEGX1_26/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2017 gnd INVX4_0/Y DFFNEGX1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2018 DFFNEGX1_26/a_66_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2019 INVX2_40/A DFFNEGX1_26/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2020 DFFNEGX1_26/a_23_6# INVX4_0/Y DFFNEGX1_26/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2021 DFFNEGX1_26/a_23_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2022 gnd DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2023 vdd DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2024 DFFNEGX1_26/a_61_74# DFFNEGX1_26/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2025 DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2026 DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2027 vdd INVX2_40/A DFFNEGX1_26/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2028 gnd INVX2_40/A DFFNEGX1_26/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2029 DFFNEGX1_26/a_61_6# DFFNEGX1_26/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2030 DFFNEGX1_26/a_76_84# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2031 INVX2_40/A DFFNEGX1_26/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2032 vdd INVX4_0/Y DFFNEGX1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2033 DFFNEGX1_26/a_31_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2034 DFFNEGX1_26/a_66_6# INVX4_0/Y DFFNEGX1_26/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2035 DFFNEGX1_26/a_17_74# OAI22X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2036 DFFNEGX1_26/a_31_74# INVX4_0/Y DFFNEGX1_26/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2037 DFFNEGX1_26/a_17_6# OAI22X1_5/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2038 INVX4_0/Y INVX4_0/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M2039 vdd INVX4_0/A INVX4_0/Y vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M2040 INVX4_0/Y INVX4_0/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M2041 gnd INVX4_0/A INVX4_0/Y Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M2042 AND2X2_2/B NAND3X1_3/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2043 NAND3X1_3/a_9_6# NAND3X1_3/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2044 AND2X2_2/B NOR2X1_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2045 AND2X2_2/B NOR2X1_10/Y NAND3X1_3/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2046 vdd NAND3X1_3/B AND2X2_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2047 NAND3X1_3/a_14_6# NAND3X1_3/B NAND3X1_3/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2048 gnd NOR2X1_28/Y AOI22X1_8/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2049 AOI22X1_8/Y NOR2X1_29/Y AOI22X1_8/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2050 AOI22X1_8/a_11_6# NOR2X1_30/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2051 AOI22X1_8/a_2_54# NOR2X1_29/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2052 AOI22X1_8/a_28_6# NOR2X1_27/Y AOI22X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2053 vdd NOR2X1_30/Y AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2054 AOI22X1_8/Y NOR2X1_27/Y AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2055 AOI22X1_8/a_2_54# NOR2X1_28/Y AOI22X1_8/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2056 OAI21X1_19/B XNOR2X1_56/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2057 NAND2X1_18/a_9_6# XNOR2X1_56/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2058 vdd XNOR2X1_55/Y OAI21X1_19/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2059 OAI21X1_19/B XNOR2X1_55/Y NAND2X1_18/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2060 gnd XNOR2X1_71/A XNOR2X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2061 out_Anum[1] XNOR2X1_71/A XNOR2X1_71/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2062 XNOR2X1_71/a_12_41# NAND3X1_8/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2063 XNOR2X1_71/a_18_54# XNOR2X1_71/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2064 XNOR2X1_71/a_35_6# XNOR2X1_71/a_2_6# out_Anum[1] Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2065 XNOR2X1_71/a_18_6# XNOR2X1_71/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2066 vdd XNOR2X1_71/A XNOR2X1_71/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2067 vdd NAND3X1_8/B XNOR2X1_71/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2068 out_Anum[1] XNOR2X1_71/a_2_6# XNOR2X1_71/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2069 XNOR2X1_71/a_35_54# XNOR2X1_71/A out_Anum[1] vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2070 XNOR2X1_71/a_12_41# NAND3X1_8/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2071 gnd NAND3X1_8/B XNOR2X1_71/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2072 gnd INVX2_54/Y XNOR2X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2073 NOR2X1_27/A INVX2_54/Y XNOR2X1_60/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2074 XNOR2X1_60/a_12_41# INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2075 XNOR2X1_60/a_18_54# XNOR2X1_60/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2076 XNOR2X1_60/a_35_6# XNOR2X1_60/a_2_6# NOR2X1_27/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2077 XNOR2X1_60/a_18_6# XNOR2X1_60/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2078 vdd INVX2_54/Y XNOR2X1_60/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2079 vdd INVX2_24/A XNOR2X1_60/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2080 NOR2X1_27/A XNOR2X1_60/a_2_6# XNOR2X1_60/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2081 XNOR2X1_60/a_35_54# INVX2_54/Y NOR2X1_27/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2082 XNOR2X1_60/a_12_41# INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2083 gnd INVX2_24/A XNOR2X1_60/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2084 gnd INVX2_56/A XNOR2X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2085 XNOR2X1_82/Y INVX2_56/A XNOR2X1_82/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2086 XNOR2X1_82/a_12_41# INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2087 XNOR2X1_82/a_18_54# XNOR2X1_82/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2088 XNOR2X1_82/a_35_6# XNOR2X1_82/a_2_6# XNOR2X1_82/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2089 XNOR2X1_82/a_18_6# XNOR2X1_82/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2090 vdd INVX2_56/A XNOR2X1_82/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2091 vdd INVX2_28/A XNOR2X1_82/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2092 XNOR2X1_82/Y XNOR2X1_82/a_2_6# XNOR2X1_82/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2093 XNOR2X1_82/a_35_54# INVX2_56/A XNOR2X1_82/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2094 XNOR2X1_82/a_12_41# INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2095 gnd INVX2_28/A XNOR2X1_82/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2096 gnd NOR2X1_0/Y OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2097 vdd OAI21X1_0/C OAI21X1_0/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2098 OAI21X1_0/Y OAI21X1_0/C OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2099 OAI21X1_0/Y INVX2_11/A OAI21X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2100 OAI21X1_0/a_9_54# NOR2X1_0/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2101 OAI21X1_0/a_2_6# INVX2_11/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2102 gnd XOR2X1_4/Y XOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2103 out_Bnum[0] XOR2X1_3/a_2_6# XOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2104 XOR2X1_3/a_13_43# XOR2X1_3/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2105 XOR2X1_3/a_18_54# XOR2X1_3/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2106 XOR2X1_3/a_35_6# XOR2X1_4/Y out_Bnum[0] Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2107 XOR2X1_3/a_18_6# XOR2X1_3/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2108 vdd XOR2X1_4/Y XOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2109 vdd XOR2X1_3/B XOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2110 out_Bnum[0] XOR2X1_4/Y XOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2111 XOR2X1_3/a_35_54# XOR2X1_3/a_2_6# out_Bnum[0] vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2112 XOR2X1_3/a_13_43# XOR2X1_3/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2113 gnd XOR2X1_3/B XOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2114 gnd MUX2X1_4/A MUX2X1_4/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2115 MUX2X1_4/a_17_50# INVX2_2/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2116 MUX2X1_4/Y MUX2X1_7/S MUX2X1_4/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2117 MUX2X1_4/a_30_54# MUX2X1_4/a_2_10# MUX2X1_4/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2118 MUX2X1_4/a_17_10# INVX2_2/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2119 vdd MUX2X1_7/S MUX2X1_4/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2120 MUX2X1_4/a_30_10# MUX2X1_7/S MUX2X1_4/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2121 gnd MUX2X1_7/S MUX2X1_4/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2122 vdd MUX2X1_4/A MUX2X1_4/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2123 MUX2X1_4/Y MUX2X1_4/a_2_10# MUX2X1_4/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2124 DFFNEGX1_16/a_76_6# INVX2_102/Y DFFNEGX1_16/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2125 gnd INVX2_102/Y DFFNEGX1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2126 DFFNEGX1_16/a_66_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2127 INVX2_30/A DFFNEGX1_16/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2128 DFFNEGX1_16/a_23_6# INVX2_102/Y DFFNEGX1_16/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2129 DFFNEGX1_16/a_23_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2130 gnd DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2131 vdd DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2132 DFFNEGX1_16/a_61_74# DFFNEGX1_16/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2133 DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2134 DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2135 vdd INVX2_30/A DFFNEGX1_16/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2136 gnd INVX2_30/A DFFNEGX1_16/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2137 DFFNEGX1_16/a_61_6# DFFNEGX1_16/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2138 DFFNEGX1_16/a_76_84# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2139 INVX2_30/A DFFNEGX1_16/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2140 vdd INVX2_102/Y DFFNEGX1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2141 DFFNEGX1_16/a_31_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2142 DFFNEGX1_16/a_66_6# INVX2_102/Y DFFNEGX1_16/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2143 DFFNEGX1_16/a_17_74# OAI22X1_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2144 DFFNEGX1_16/a_31_74# INVX2_102/Y DFFNEGX1_16/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2145 DFFNEGX1_16/a_17_6# OAI22X1_11/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2146 DFFNEGX1_38/a_76_6# INVX4_0/Y DFFNEGX1_38/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2147 gnd INVX4_0/Y DFFNEGX1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2148 DFFNEGX1_38/a_66_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2149 INVX2_55/A DFFNEGX1_38/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2150 DFFNEGX1_38/a_23_6# INVX4_0/Y DFFNEGX1_38/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2151 DFFNEGX1_38/a_23_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2152 gnd DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2153 vdd DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2154 DFFNEGX1_38/a_61_74# DFFNEGX1_38/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2155 DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2156 DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2157 vdd INVX2_55/A DFFNEGX1_38/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2158 gnd INVX2_55/A DFFNEGX1_38/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2159 DFFNEGX1_38/a_61_6# DFFNEGX1_38/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2160 DFFNEGX1_38/a_76_84# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2161 INVX2_55/A DFFNEGX1_38/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2162 vdd INVX4_0/Y DFFNEGX1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2163 DFFNEGX1_38/a_31_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2164 DFFNEGX1_38/a_66_6# INVX4_0/Y DFFNEGX1_38/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2165 DFFNEGX1_38/a_17_74# OAI22X1_25/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2166 DFFNEGX1_38/a_31_74# INVX4_0/Y DFFNEGX1_38/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2167 DFFNEGX1_38/a_17_6# OAI22X1_25/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2168 DFFNEGX1_27/a_76_6# INVX4_0/Y DFFNEGX1_27/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2169 gnd INVX4_0/Y DFFNEGX1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2170 DFFNEGX1_27/a_66_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2171 INVX2_41/A DFFNEGX1_27/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2172 DFFNEGX1_27/a_23_6# INVX4_0/Y DFFNEGX1_27/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2173 DFFNEGX1_27/a_23_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2174 gnd DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2175 vdd DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2176 DFFNEGX1_27/a_61_74# DFFNEGX1_27/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2177 DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2178 DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2179 vdd INVX2_41/A DFFNEGX1_27/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2180 gnd INVX2_41/A DFFNEGX1_27/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2181 DFFNEGX1_27/a_61_6# DFFNEGX1_27/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2182 DFFNEGX1_27/a_76_84# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2183 INVX2_41/A DFFNEGX1_27/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2184 vdd INVX4_0/Y DFFNEGX1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2185 DFFNEGX1_27/a_31_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2186 DFFNEGX1_27/a_66_6# INVX4_0/Y DFFNEGX1_27/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2187 DFFNEGX1_27/a_17_74# OAI22X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2188 DFFNEGX1_27/a_31_74# INVX4_0/Y DFFNEGX1_27/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2189 DFFNEGX1_27/a_17_6# OAI22X1_4/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2190 OAI21X1_5/A INVX2_21/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2191 NAND3X1_4/a_9_6# INVX2_21/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2192 OAI21X1_5/A AND2X2_3/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2193 OAI21X1_5/A AND2X2_3/Y NAND3X1_4/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2194 vdd INVX2_70/A OAI21X1_5/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2195 NAND3X1_4/a_14_6# INVX2_70/A NAND3X1_4/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2196 OAI21X1_19/A XNOR2X1_58/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2197 NAND2X1_19/a_9_6# XNOR2X1_58/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2198 vdd XNOR2X1_57/Y OAI21X1_19/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2199 OAI21X1_19/A XNOR2X1_57/Y NAND2X1_19/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2200 gnd INVX2_47/Y XNOR2X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2201 NOR2X1_33/B INVX2_47/Y XNOR2X1_83/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2202 XNOR2X1_83/a_12_41# INVX2_23/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2203 XNOR2X1_83/a_18_54# XNOR2X1_83/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2204 XNOR2X1_83/a_35_6# XNOR2X1_83/a_2_6# NOR2X1_33/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2205 XNOR2X1_83/a_18_6# XNOR2X1_83/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2206 vdd INVX2_47/Y XNOR2X1_83/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2207 vdd INVX2_23/A XNOR2X1_83/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2208 NOR2X1_33/B XNOR2X1_83/a_2_6# XNOR2X1_83/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2209 XNOR2X1_83/a_35_54# INVX2_47/Y NOR2X1_33/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2210 XNOR2X1_83/a_12_41# INVX2_23/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2211 gnd INVX2_23/A XNOR2X1_83/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2212 gnd INVX2_56/Y XNOR2X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2213 NOR2X1_28/B INVX2_56/Y XNOR2X1_61/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2214 XNOR2X1_61/a_12_41# INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2215 XNOR2X1_61/a_18_54# XNOR2X1_61/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2216 XNOR2X1_61/a_35_6# XNOR2X1_61/a_2_6# NOR2X1_28/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2217 XNOR2X1_61/a_18_6# XNOR2X1_61/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2218 vdd INVX2_56/Y XNOR2X1_61/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2219 vdd INVX2_26/A XNOR2X1_61/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2220 NOR2X1_28/B XNOR2X1_61/a_2_6# XNOR2X1_61/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2221 XNOR2X1_61/a_35_54# INVX2_56/Y NOR2X1_28/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2222 XNOR2X1_61/a_12_41# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2223 gnd INVX2_26/A XNOR2X1_61/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2224 gnd INVX2_43/A XNOR2X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2225 out_Anum[0] INVX2_43/A XNOR2X1_72/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2226 XNOR2X1_72/a_12_41# NAND3X1_8/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2227 XNOR2X1_72/a_18_54# XNOR2X1_72/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2228 XNOR2X1_72/a_35_6# XNOR2X1_72/a_2_6# out_Anum[0] Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2229 XNOR2X1_72/a_18_6# XNOR2X1_72/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2230 vdd INVX2_43/A XNOR2X1_72/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2231 vdd NAND3X1_8/A XNOR2X1_72/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2232 out_Anum[0] XNOR2X1_72/a_2_6# XNOR2X1_72/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2233 XNOR2X1_72/a_35_54# INVX2_43/A out_Anum[0] vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2234 XNOR2X1_72/a_12_41# NAND3X1_8/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2235 gnd NAND3X1_8/A XNOR2X1_72/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2236 gnd INVX2_55/Y XNOR2X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2237 NOR2X1_24/A INVX2_55/Y XNOR2X1_50/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2238 XNOR2X1_50/a_12_41# INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2239 XNOR2X1_50/a_18_54# XNOR2X1_50/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2240 XNOR2X1_50/a_35_6# XNOR2X1_50/a_2_6# NOR2X1_24/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2241 XNOR2X1_50/a_18_6# XNOR2X1_50/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2242 vdd INVX2_55/Y XNOR2X1_50/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2243 vdd INVX2_32/A XNOR2X1_50/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2244 NOR2X1_24/A XNOR2X1_50/a_2_6# XNOR2X1_50/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2245 XNOR2X1_50/a_35_54# INVX2_55/Y NOR2X1_24/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2246 XNOR2X1_50/a_12_41# INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2247 gnd INVX2_32/A XNOR2X1_50/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2248 gnd NOR2X1_1/Y OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2249 vdd MUX2X1_8/Y OAI21X1_1/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2250 OAI21X1_1/Y MUX2X1_8/Y OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2251 OAI21X1_1/Y INVX2_8/A OAI21X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2252 OAI21X1_1/a_9_54# NOR2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2253 OAI21X1_1/a_2_6# INVX2_8/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2254 gnd MUX2X1_5/A MUX2X1_5/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2255 MUX2X1_5/a_17_50# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2256 INVX2_5/A MUX2X1_7/S MUX2X1_5/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2257 MUX2X1_5/a_30_54# MUX2X1_5/a_2_10# INVX2_5/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2258 MUX2X1_5/a_17_10# INVX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2259 vdd MUX2X1_7/S MUX2X1_5/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2260 MUX2X1_5/a_30_10# MUX2X1_7/S INVX2_5/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2261 gnd MUX2X1_7/S MUX2X1_5/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2262 vdd MUX2X1_5/A MUX2X1_5/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2263 INVX2_5/A MUX2X1_5/a_2_10# MUX2X1_5/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2264 gnd XOR2X1_4/A XOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2265 XOR2X1_4/Y XOR2X1_4/a_2_6# XOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2266 XOR2X1_4/a_13_43# XOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2267 XOR2X1_4/a_18_54# XOR2X1_4/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2268 XOR2X1_4/a_35_6# XOR2X1_4/A XOR2X1_4/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2269 XOR2X1_4/a_18_6# XOR2X1_4/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2270 vdd XOR2X1_4/A XOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2271 vdd XOR2X1_5/Y XOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2272 XOR2X1_4/Y XOR2X1_4/A XOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2273 XOR2X1_4/a_35_54# XOR2X1_4/a_2_6# XOR2X1_4/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2274 XOR2X1_4/a_13_43# XOR2X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2275 gnd XOR2X1_5/Y XOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2276 OAI22X1_6/A AND2X2_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2277 OAI22X1_6/A AND2X2_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2278 DFFNEGX1_39/a_76_6# INVX4_0/Y DFFNEGX1_39/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2279 gnd INVX4_0/Y DFFNEGX1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2280 DFFNEGX1_39/a_66_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2281 INVX2_56/A DFFNEGX1_39/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2282 DFFNEGX1_39/a_23_6# INVX4_0/Y DFFNEGX1_39/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2283 DFFNEGX1_39/a_23_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2284 gnd DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2285 vdd DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2286 DFFNEGX1_39/a_61_74# DFFNEGX1_39/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2287 DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2288 DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2289 vdd INVX2_56/A DFFNEGX1_39/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2290 gnd INVX2_56/A DFFNEGX1_39/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2291 DFFNEGX1_39/a_61_6# DFFNEGX1_39/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2292 DFFNEGX1_39/a_76_84# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2293 INVX2_56/A DFFNEGX1_39/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2294 vdd INVX4_0/Y DFFNEGX1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2295 DFFNEGX1_39/a_31_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2296 DFFNEGX1_39/a_66_6# INVX4_0/Y DFFNEGX1_39/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2297 DFFNEGX1_39/a_17_74# OAI22X1_24/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2298 DFFNEGX1_39/a_31_74# INVX4_0/Y DFFNEGX1_39/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2299 DFFNEGX1_39/a_17_6# OAI22X1_24/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2300 DFFNEGX1_17/a_76_6# INVX2_102/Y DFFNEGX1_17/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2301 gnd INVX2_102/Y DFFNEGX1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2302 DFFNEGX1_17/a_66_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2303 INVX2_31/A DFFNEGX1_17/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2304 DFFNEGX1_17/a_23_6# INVX2_102/Y DFFNEGX1_17/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2305 DFFNEGX1_17/a_23_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2306 gnd DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2307 vdd DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2308 DFFNEGX1_17/a_61_74# DFFNEGX1_17/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2309 DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2310 DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2311 vdd INVX2_31/A DFFNEGX1_17/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2312 gnd INVX2_31/A DFFNEGX1_17/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2313 DFFNEGX1_17/a_61_6# DFFNEGX1_17/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2314 DFFNEGX1_17/a_76_84# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2315 INVX2_31/A DFFNEGX1_17/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2316 vdd INVX2_102/Y DFFNEGX1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2317 DFFNEGX1_17/a_31_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2318 DFFNEGX1_17/a_66_6# INVX2_102/Y DFFNEGX1_17/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2319 DFFNEGX1_17/a_17_74# OAI22X1_17/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2320 DFFNEGX1_17/a_31_74# INVX2_102/Y DFFNEGX1_17/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2321 DFFNEGX1_17/a_17_6# OAI22X1_17/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2322 DFFNEGX1_28/a_76_6# INVX4_0/Y DFFNEGX1_28/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2323 gnd INVX4_0/Y DFFNEGX1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2324 DFFNEGX1_28/a_66_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2325 INVX2_42/A DFFNEGX1_28/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2326 DFFNEGX1_28/a_23_6# INVX4_0/Y DFFNEGX1_28/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2327 DFFNEGX1_28/a_23_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2328 gnd DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2329 vdd DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2330 DFFNEGX1_28/a_61_74# DFFNEGX1_28/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2331 DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2332 DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2333 vdd INVX2_42/A DFFNEGX1_28/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2334 gnd INVX2_42/A DFFNEGX1_28/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2335 DFFNEGX1_28/a_61_6# DFFNEGX1_28/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2336 DFFNEGX1_28/a_76_84# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2337 INVX2_42/A DFFNEGX1_28/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2338 vdd INVX4_0/Y DFFNEGX1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2339 DFFNEGX1_28/a_31_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2340 DFFNEGX1_28/a_66_6# INVX4_0/Y DFFNEGX1_28/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2341 DFFNEGX1_28/a_17_74# OAI22X1_3/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2342 DFFNEGX1_28/a_31_74# INVX4_0/Y DFFNEGX1_28/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2343 DFFNEGX1_28/a_17_6# OAI22X1_3/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2344 AND2X2_3/B NAND3X1_5/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2345 NAND3X1_5/a_9_6# NAND3X1_5/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2346 AND2X2_3/B NOR2X1_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2347 AND2X2_3/B NOR2X1_11/Y NAND3X1_5/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2348 vdd NAND3X1_5/B AND2X2_3/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2349 NAND3X1_5/a_14_6# NAND3X1_5/B NAND3X1_5/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2350 gnd INVX2_44/Y XNOR2X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2351 NOR2X1_33/A INVX2_44/Y XNOR2X1_84/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2352 XNOR2X1_84/a_12_41# INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2353 XNOR2X1_84/a_18_54# XNOR2X1_84/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2354 XNOR2X1_84/a_35_6# XNOR2X1_84/a_2_6# NOR2X1_33/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2355 XNOR2X1_84/a_18_6# XNOR2X1_84/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2356 vdd INVX2_44/Y XNOR2X1_84/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2357 vdd INVX2_24/A XNOR2X1_84/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2358 NOR2X1_33/A XNOR2X1_84/a_2_6# XNOR2X1_84/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2359 XNOR2X1_84/a_35_54# INVX2_44/Y NOR2X1_33/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2360 XNOR2X1_84/a_12_41# INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2361 gnd INVX2_24/A XNOR2X1_84/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2362 gnd INVX2_48/Y XNOR2X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2363 NAND3X1_8/A INVX2_48/Y XNOR2X1_73/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2364 XNOR2X1_73/a_12_41# XNOR2X1_74/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2365 XNOR2X1_73/a_18_54# XNOR2X1_73/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2366 XNOR2X1_73/a_35_6# XNOR2X1_73/a_2_6# NAND3X1_8/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2367 XNOR2X1_73/a_18_6# XNOR2X1_73/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2368 vdd INVX2_48/Y XNOR2X1_73/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2369 vdd XNOR2X1_74/Y XNOR2X1_73/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2370 NAND3X1_8/A XNOR2X1_73/a_2_6# XNOR2X1_73/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2371 XNOR2X1_73/a_35_54# INVX2_48/Y NAND3X1_8/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2372 XNOR2X1_73/a_12_41# XNOR2X1_74/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2373 gnd XNOR2X1_74/Y XNOR2X1_73/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2374 gnd INVX2_39/Y XNOR2X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2375 NOR2X1_21/A INVX2_39/Y XNOR2X1_40/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2376 XNOR2X1_40/a_12_41# INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2377 XNOR2X1_40/a_18_54# XNOR2X1_40/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2378 XNOR2X1_40/a_35_6# XNOR2X1_40/a_2_6# NOR2X1_21/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2379 XNOR2X1_40/a_18_6# XNOR2X1_40/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2380 vdd INVX2_39/Y XNOR2X1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2381 vdd INVX2_30/A XNOR2X1_40/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2382 NOR2X1_21/A XNOR2X1_40/a_2_6# XNOR2X1_40/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2383 XNOR2X1_40/a_35_54# INVX2_39/Y NOR2X1_21/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2384 XNOR2X1_40/a_12_41# INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2385 gnd INVX2_30/A XNOR2X1_40/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2386 gnd INVX2_55/Y XNOR2X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2387 NOR2X1_28/A INVX2_55/Y XNOR2X1_62/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2388 XNOR2X1_62/a_12_41# INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2389 XNOR2X1_62/a_18_54# XNOR2X1_62/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2390 XNOR2X1_62/a_35_6# XNOR2X1_62/a_2_6# NOR2X1_28/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2391 XNOR2X1_62/a_18_6# XNOR2X1_62/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2392 vdd INVX2_55/Y XNOR2X1_62/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2393 vdd INVX2_25/A XNOR2X1_62/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2394 NOR2X1_28/A XNOR2X1_62/a_2_6# XNOR2X1_62/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2395 XNOR2X1_62/a_35_54# INVX2_55/Y NOR2X1_28/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2396 XNOR2X1_62/a_12_41# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2397 gnd INVX2_25/A XNOR2X1_62/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2398 gnd INVX2_42/Y XNOR2X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2399 NOR2X1_25/B INVX2_42/Y XNOR2X1_51/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2400 XNOR2X1_51/a_12_41# INVX2_18/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2401 XNOR2X1_51/a_18_54# XNOR2X1_51/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2402 XNOR2X1_51/a_35_6# XNOR2X1_51/a_2_6# NOR2X1_25/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2403 XNOR2X1_51/a_18_6# XNOR2X1_51/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2404 vdd INVX2_42/Y XNOR2X1_51/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2405 vdd INVX2_18/A XNOR2X1_51/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2406 NOR2X1_25/B XNOR2X1_51/a_2_6# XNOR2X1_51/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2407 XNOR2X1_51/a_35_54# INVX2_42/Y NOR2X1_25/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2408 XNOR2X1_51/a_12_41# INVX2_18/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2409 gnd INVX2_18/A XNOR2X1_51/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2410 gnd NOR2X1_2/Y OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2411 vdd MUX2X1_4/Y MUX2X1_9/S vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2412 MUX2X1_9/S MUX2X1_4/Y OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2413 MUX2X1_9/S INVX2_5/A OAI21X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2414 OAI21X1_2/a_9_54# NOR2X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2415 OAI21X1_2/a_2_6# INVX2_5/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2416 DFFNEGX1_0/a_76_6# INVX2_101/Y DFFNEGX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2417 gnd INVX2_101/Y DFFNEGX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2418 DFFNEGX1_0/a_66_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2419 AOI22X1_3/C DFFNEGX1_0/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2420 DFFNEGX1_0/a_23_6# INVX2_101/Y DFFNEGX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2421 DFFNEGX1_0/a_23_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2422 gnd DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2423 vdd DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2424 DFFNEGX1_0/a_61_74# DFFNEGX1_0/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2425 DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2426 DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2427 vdd AOI22X1_3/C DFFNEGX1_0/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2428 gnd AOI22X1_3/C DFFNEGX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2429 DFFNEGX1_0/a_61_6# DFFNEGX1_0/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2430 DFFNEGX1_0/a_76_84# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2431 AOI22X1_3/C DFFNEGX1_0/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2432 vdd INVX2_101/Y DFFNEGX1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2433 DFFNEGX1_0/a_31_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2434 DFFNEGX1_0/a_66_6# INVX2_101/Y DFFNEGX1_0/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2435 DFFNEGX1_0/a_17_74# INVX2_77/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2436 DFFNEGX1_0/a_31_74# INVX2_101/Y DFFNEGX1_0/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2437 DFFNEGX1_0/a_17_6# INVX2_77/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2438 gnd XOR2X1_5/A XOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2439 XOR2X1_5/Y XOR2X1_5/a_2_6# XOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2440 XOR2X1_5/a_13_43# XOR2X1_5/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2441 XOR2X1_5/a_18_54# XOR2X1_5/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2442 XOR2X1_5/a_35_6# XOR2X1_5/A XOR2X1_5/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2443 XOR2X1_5/a_18_6# XOR2X1_5/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2444 vdd XOR2X1_5/A XOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2445 vdd XOR2X1_5/B XOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2446 XOR2X1_5/Y XOR2X1_5/A XOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2447 XOR2X1_5/a_35_54# XOR2X1_5/a_2_6# XOR2X1_5/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2448 XOR2X1_5/a_13_43# XOR2X1_5/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2449 gnd XOR2X1_5/B XOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2450 gnd INVX2_4/A MUX2X1_6/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2451 MUX2X1_6/a_17_50# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2452 INVX2_6/A MUX2X1_7/S MUX2X1_6/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2453 MUX2X1_6/a_30_54# MUX2X1_6/a_2_10# INVX2_6/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2454 MUX2X1_6/a_17_10# INVX2_4/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2455 vdd MUX2X1_7/S MUX2X1_6/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2456 MUX2X1_6/a_30_10# MUX2X1_7/S INVX2_6/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2457 gnd MUX2X1_7/S MUX2X1_6/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2458 vdd INVX2_4/A MUX2X1_6/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2459 INVX2_6/A MUX2X1_6/a_2_10# MUX2X1_6/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2460 INVX2_101/Y BUFX2_1/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2461 INVX2_101/Y BUFX2_1/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2462 DFFNEGX1_18/a_76_6# INVX2_102/Y DFFNEGX1_18/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2463 gnd INVX2_102/Y DFFNEGX1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2464 DFFNEGX1_18/a_66_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2465 INVX2_32/A DFFNEGX1_18/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2466 DFFNEGX1_18/a_23_6# INVX2_102/Y DFFNEGX1_18/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2467 DFFNEGX1_18/a_23_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2468 gnd DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2469 vdd DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2470 DFFNEGX1_18/a_61_74# DFFNEGX1_18/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2471 DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2472 DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2473 vdd INVX2_32/A DFFNEGX1_18/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2474 gnd INVX2_32/A DFFNEGX1_18/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2475 DFFNEGX1_18/a_61_6# DFFNEGX1_18/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2476 DFFNEGX1_18/a_76_84# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2477 INVX2_32/A DFFNEGX1_18/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2478 vdd INVX2_102/Y DFFNEGX1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2479 DFFNEGX1_18/a_31_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2480 DFFNEGX1_18/a_66_6# INVX2_102/Y DFFNEGX1_18/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2481 DFFNEGX1_18/a_17_74# OAI22X1_16/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2482 DFFNEGX1_18/a_31_74# INVX2_102/Y DFFNEGX1_18/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2483 DFFNEGX1_18/a_17_6# OAI22X1_16/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2484 DFFNEGX1_29/a_76_6# INVX4_0/Y DFFNEGX1_29/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2485 gnd INVX4_0/Y DFFNEGX1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2486 DFFNEGX1_29/a_66_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2487 INVX2_44/A DFFNEGX1_29/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2488 DFFNEGX1_29/a_23_6# INVX4_0/Y DFFNEGX1_29/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2489 DFFNEGX1_29/a_23_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2490 gnd DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2491 vdd DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2492 DFFNEGX1_29/a_61_74# DFFNEGX1_29/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2493 DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2494 DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2495 vdd INVX2_44/A DFFNEGX1_29/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2496 gnd INVX2_44/A DFFNEGX1_29/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2497 DFFNEGX1_29/a_61_6# DFFNEGX1_29/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2498 DFFNEGX1_29/a_76_84# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2499 INVX2_44/A DFFNEGX1_29/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2500 vdd INVX4_0/Y DFFNEGX1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2501 DFFNEGX1_29/a_31_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2502 DFFNEGX1_29/a_66_6# INVX4_0/Y DFFNEGX1_29/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2503 DFFNEGX1_29/a_17_74# OAI22X1_2/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2504 DFFNEGX1_29/a_31_74# INVX4_0/Y DFFNEGX1_29/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2505 DFFNEGX1_29/a_17_6# OAI22X1_2/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2506 INVX2_97/A NOR2X1_9/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2507 NAND3X1_6/a_9_6# NOR2X1_9/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2508 INVX2_97/A NOR2X1_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2509 INVX2_97/A NOR2X1_13/Y NAND3X1_6/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2510 vdd NOR2X1_14/Y INVX2_97/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2511 NAND3X1_6/a_14_6# NOR2X1_14/Y NAND3X1_6/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2512 vdd BUFX2_1/A BUFX2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0.11n pd=46u as=100p ps=50u
M2513 gnd BUFX2_1/A BUFX2_0/a_2_6# Gnd nfet w=10 l=2
+  ad=55p pd=26u as=50p ps=30u
M2514 BUFX2_0/Y BUFX2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.11n ps=46u
M2515 BUFX2_0/Y BUFX2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=55p ps=26u
M2516 AOI21X1_0/a_2_54# INVX2_72/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M2517 AOI21X1_0/a_12_6# NOR2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M2518 gnd INVX2_73/A NOR2X1_6/A Gnd nfet w=10 l=2
+  ad=50p pd=30u as=55p ps=26u
M2519 vdd NOR2X1_7/A AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M2520 NOR2X1_6/A INVX2_73/A AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M2521 NOR2X1_6/A INVX2_72/Y AOI21X1_0/a_12_6# Gnd nfet w=20 l=2
+  ad=55p pd=26u as=29.999998p ps=23u
M2522 INVX2_0/Y INVX2_0/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2523 INVX2_0/Y INVX2_0/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2524 gnd INVX2_55/Y XNOR2X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2525 NOR2X1_18/A INVX2_55/Y XNOR2X1_30/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2526 XNOR2X1_30/a_12_41# INVX2_36/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2527 XNOR2X1_30/a_18_54# XNOR2X1_30/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2528 XNOR2X1_30/a_35_6# XNOR2X1_30/a_2_6# NOR2X1_18/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2529 XNOR2X1_30/a_18_6# XNOR2X1_30/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2530 vdd INVX2_55/Y XNOR2X1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2531 vdd INVX2_36/A XNOR2X1_30/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2532 NOR2X1_18/A XNOR2X1_30/a_2_6# XNOR2X1_30/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2533 XNOR2X1_30/a_35_54# INVX2_55/Y NOR2X1_18/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2534 XNOR2X1_30/a_12_41# INVX2_36/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2535 gnd INVX2_36/A XNOR2X1_30/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2536 gnd INVX2_41/Y XNOR2X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2537 NOR2X1_22/B INVX2_41/Y XNOR2X1_41/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2538 XNOR2X1_41/a_12_41# INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2539 XNOR2X1_41/a_18_54# XNOR2X1_41/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2540 XNOR2X1_41/a_35_6# XNOR2X1_41/a_2_6# NOR2X1_22/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2541 XNOR2X1_41/a_18_6# XNOR2X1_41/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2542 vdd INVX2_41/Y XNOR2X1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2543 vdd INVX2_28/A XNOR2X1_41/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2544 NOR2X1_22/B XNOR2X1_41/a_2_6# XNOR2X1_41/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2545 XNOR2X1_41/a_35_54# INVX2_41/Y NOR2X1_22/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2546 XNOR2X1_41/a_12_41# INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2547 gnd INVX2_28/A XNOR2X1_41/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2548 gnd INVX2_60/Y XNOR2X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2549 XNOR2X1_74/Y INVX2_60/Y XNOR2X1_74/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2550 XNOR2X1_74/a_12_41# INVX2_53/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2551 XNOR2X1_74/a_18_54# XNOR2X1_74/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2552 XNOR2X1_74/a_35_6# XNOR2X1_74/a_2_6# XNOR2X1_74/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2553 XNOR2X1_74/a_18_6# XNOR2X1_74/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2554 vdd INVX2_60/Y XNOR2X1_74/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2555 vdd INVX2_53/Y XNOR2X1_74/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2556 XNOR2X1_74/Y XNOR2X1_74/a_2_6# XNOR2X1_74/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2557 XNOR2X1_74/a_35_54# INVX2_60/Y XNOR2X1_74/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2558 XNOR2X1_74/a_12_41# INVX2_53/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2559 gnd INVX2_53/Y XNOR2X1_74/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2560 gnd INVX2_45/A XNOR2X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2561 XNOR2X1_85/Y INVX2_45/A XNOR2X1_85/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2562 XNOR2X1_85/a_12_41# INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2563 XNOR2X1_85/a_18_54# XNOR2X1_85/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2564 XNOR2X1_85/a_35_6# XNOR2X1_85/a_2_6# XNOR2X1_85/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2565 XNOR2X1_85/a_18_6# XNOR2X1_85/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2566 vdd INVX2_45/A XNOR2X1_85/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2567 vdd INVX2_25/A XNOR2X1_85/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2568 XNOR2X1_85/Y XNOR2X1_85/a_2_6# XNOR2X1_85/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2569 XNOR2X1_85/a_35_54# INVX2_45/A XNOR2X1_85/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2570 XNOR2X1_85/a_12_41# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2571 gnd INVX2_25/A XNOR2X1_85/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2572 gnd INVX2_42/Y XNOR2X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2573 NOR2X1_29/B INVX2_42/Y XNOR2X1_63/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2574 XNOR2X1_63/a_12_41# INVX2_23/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2575 XNOR2X1_63/a_18_54# XNOR2X1_63/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2576 XNOR2X1_63/a_35_6# XNOR2X1_63/a_2_6# NOR2X1_29/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2577 XNOR2X1_63/a_18_6# XNOR2X1_63/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2578 vdd INVX2_42/Y XNOR2X1_63/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2579 vdd INVX2_23/A XNOR2X1_63/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2580 NOR2X1_29/B XNOR2X1_63/a_2_6# XNOR2X1_63/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2581 XNOR2X1_63/a_35_54# INVX2_42/Y NOR2X1_29/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2582 XNOR2X1_63/a_12_41# INVX2_23/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2583 gnd INVX2_23/A XNOR2X1_63/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2584 gnd INVX2_39/Y XNOR2X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2585 NOR2X1_25/A INVX2_39/Y XNOR2X1_52/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2586 XNOR2X1_52/a_12_41# INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2587 XNOR2X1_52/a_18_54# XNOR2X1_52/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2588 XNOR2X1_52/a_35_6# XNOR2X1_52/a_2_6# NOR2X1_25/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2589 XNOR2X1_52/a_18_6# XNOR2X1_52/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2590 vdd INVX2_39/Y XNOR2X1_52/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2591 vdd INVX2_33/A XNOR2X1_52/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2592 NOR2X1_25/A XNOR2X1_52/a_2_6# XNOR2X1_52/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2593 XNOR2X1_52/a_35_54# INVX2_39/Y NOR2X1_25/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2594 XNOR2X1_52/a_12_41# INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2595 gnd INVX2_33/A XNOR2X1_52/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2596 gnd NOR2X1_3/Y OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2597 vdd MUX2X1_0/Y MUX2X1_7/S vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2598 MUX2X1_7/S MUX2X1_0/Y OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2599 MUX2X1_7/S INVX2_2/A OAI21X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2600 OAI21X1_3/a_9_54# NOR2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2601 OAI21X1_3/a_2_6# INVX2_2/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2602 DFFNEGX1_1/a_76_6# INVX2_101/Y DFFNEGX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2603 gnd INVX2_101/Y DFFNEGX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2604 DFFNEGX1_1/a_66_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2605 NAND2X1_2/A DFFNEGX1_1/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2606 DFFNEGX1_1/a_23_6# INVX2_101/Y DFFNEGX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2607 DFFNEGX1_1/a_23_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2608 gnd DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2609 vdd DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2610 DFFNEGX1_1/a_61_74# DFFNEGX1_1/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2611 DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2612 DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2613 vdd NAND2X1_2/A DFFNEGX1_1/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2614 gnd NAND2X1_2/A DFFNEGX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2615 DFFNEGX1_1/a_61_6# DFFNEGX1_1/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2616 DFFNEGX1_1/a_76_84# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2617 NAND2X1_2/A DFFNEGX1_1/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2618 vdd INVX2_101/Y DFFNEGX1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2619 DFFNEGX1_1/a_31_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2620 DFFNEGX1_1/a_66_6# INVX2_101/Y DFFNEGX1_1/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2621 DFFNEGX1_1/a_17_74# INVX2_76/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2622 DFFNEGX1_1/a_31_74# INVX2_101/Y DFFNEGX1_1/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2623 DFFNEGX1_1/a_17_6# INVX2_76/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2624 gnd DFFSR_4/D MUX2X1_7/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2625 MUX2X1_7/a_17_50# DFFSR_4/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2626 INVX2_7/A MUX2X1_7/S MUX2X1_7/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2627 MUX2X1_7/a_30_54# MUX2X1_7/a_2_10# INVX2_7/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2628 MUX2X1_7/a_17_10# DFFSR_4/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2629 vdd MUX2X1_7/S MUX2X1_7/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2630 MUX2X1_7/a_30_10# MUX2X1_7/S INVX2_7/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2631 gnd MUX2X1_7/S MUX2X1_7/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2632 vdd DFFSR_4/D MUX2X1_7/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2633 INVX2_7/A MUX2X1_7/a_2_10# MUX2X1_7/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2634 INVX2_102/Y BUFX2_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2635 INVX2_102/Y BUFX2_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2636 DFFNEGX1_19/a_76_6# INVX2_102/Y DFFNEGX1_19/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2637 gnd INVX2_102/Y DFFNEGX1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2638 DFFNEGX1_19/a_66_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2639 INVX2_33/A DFFNEGX1_19/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2640 DFFNEGX1_19/a_23_6# INVX2_102/Y DFFNEGX1_19/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2641 DFFNEGX1_19/a_23_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2642 gnd DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2643 vdd DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2644 DFFNEGX1_19/a_61_74# DFFNEGX1_19/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2645 DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2646 DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2647 vdd INVX2_33/A DFFNEGX1_19/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2648 gnd INVX2_33/A DFFNEGX1_19/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2649 DFFNEGX1_19/a_61_6# DFFNEGX1_19/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2650 DFFNEGX1_19/a_76_84# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2651 INVX2_33/A DFFNEGX1_19/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2652 vdd INVX2_102/Y DFFNEGX1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2653 DFFNEGX1_19/a_31_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2654 DFFNEGX1_19/a_66_6# INVX2_102/Y DFFNEGX1_19/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2655 DFFNEGX1_19/a_17_74# OAI22X1_15/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2656 DFFNEGX1_19/a_31_74# INVX2_102/Y DFFNEGX1_19/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2657 DFFNEGX1_19/a_17_6# OAI22X1_15/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2658 INVX2_59/A XOR2X1_3/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2659 NAND3X1_7/a_9_6# XOR2X1_3/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2660 INVX2_59/A XOR2X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2661 INVX2_59/A XOR2X1_4/Y NAND3X1_7/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2662 vdd INVX2_58/Y INVX2_59/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2663 NAND3X1_7/a_14_6# INVX2_58/Y NAND3X1_7/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2664 vdd BUFX2_1/A BUFX2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2665 gnd BUFX2_1/A BUFX2_1/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2666 BUFX2_1/Y BUFX2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2667 BUFX2_1/Y BUFX2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2668 INVX2_1/Y INVX2_1/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2669 INVX2_1/Y INVX2_1/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2670 AOI21X1_1/a_2_54# NOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M2671 AOI21X1_1/a_12_6# INVX2_34/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2672 gnd OR2X1_0/Y AOI21X1_1/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M2673 vdd INVX2_34/Y AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2674 AOI21X1_1/Y OR2X1_0/Y AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2675 AOI21X1_1/Y NOR2X1_8/Y AOI21X1_1/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2676 gnd NAND2X1_3/A XNOR2X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2677 NAND3X1_5/B NAND2X1_3/A XNOR2X1_20/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2678 XNOR2X1_20/a_12_41# INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2679 XNOR2X1_20/a_18_54# XNOR2X1_20/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2680 XNOR2X1_20/a_35_6# XNOR2X1_20/a_2_6# NAND3X1_5/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2681 XNOR2X1_20/a_18_6# XNOR2X1_20/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2682 vdd NAND2X1_3/A XNOR2X1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2683 vdd INVX2_25/A XNOR2X1_20/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2684 NAND3X1_5/B XNOR2X1_20/a_2_6# XNOR2X1_20/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2685 XNOR2X1_20/a_35_54# NAND2X1_3/A NAND3X1_5/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2686 XNOR2X1_20/a_12_41# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2687 gnd INVX2_25/A XNOR2X1_20/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2688 gnd INVX2_52/Y XNOR2X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2689 NOR2X1_31/B INVX2_52/Y XNOR2X1_75/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2690 XNOR2X1_75/a_12_41# INVX2_18/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2691 XNOR2X1_75/a_18_54# XNOR2X1_75/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2692 XNOR2X1_75/a_35_6# XNOR2X1_75/a_2_6# NOR2X1_31/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2693 XNOR2X1_75/a_18_6# XNOR2X1_75/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2694 vdd INVX2_52/Y XNOR2X1_75/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2695 vdd INVX2_18/A XNOR2X1_75/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2696 NOR2X1_31/B XNOR2X1_75/a_2_6# XNOR2X1_75/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2697 XNOR2X1_75/a_35_54# INVX2_52/Y NOR2X1_31/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2698 XNOR2X1_75/a_12_41# INVX2_18/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2699 gnd INVX2_18/A XNOR2X1_75/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2700 gnd INVX2_36/A XNOR2X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2701 XNOR2X1_31/Y INVX2_36/A XNOR2X1_31/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2702 XNOR2X1_31/a_12_41# INVX2_45/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2703 XNOR2X1_31/a_18_54# XNOR2X1_31/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2704 XNOR2X1_31/a_35_6# XNOR2X1_31/a_2_6# XNOR2X1_31/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2705 XNOR2X1_31/a_18_6# XNOR2X1_31/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2706 vdd INVX2_36/A XNOR2X1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2707 vdd INVX2_45/A XNOR2X1_31/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2708 XNOR2X1_31/Y XNOR2X1_31/a_2_6# XNOR2X1_31/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2709 XNOR2X1_31/a_35_54# INVX2_36/A XNOR2X1_31/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2710 XNOR2X1_31/a_12_41# INVX2_45/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2711 gnd INVX2_45/A XNOR2X1_31/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2712 gnd INVX2_39/Y XNOR2X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2713 NOR2X1_29/A INVX2_39/Y XNOR2X1_64/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2714 XNOR2X1_64/a_12_41# INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2715 XNOR2X1_64/a_18_54# XNOR2X1_64/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2716 XNOR2X1_64/a_35_6# XNOR2X1_64/a_2_6# NOR2X1_29/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2717 XNOR2X1_64/a_18_6# XNOR2X1_64/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2718 vdd INVX2_39/Y XNOR2X1_64/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2719 vdd INVX2_24/A XNOR2X1_64/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2720 NOR2X1_29/A XNOR2X1_64/a_2_6# XNOR2X1_64/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2721 XNOR2X1_64/a_35_54# INVX2_39/Y NOR2X1_29/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2722 XNOR2X1_64/a_12_41# INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2723 gnd INVX2_24/A XNOR2X1_64/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2724 gnd INVX2_41/Y XNOR2X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2725 NOR2X1_26/B INVX2_41/Y XNOR2X1_53/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2726 XNOR2X1_53/a_12_41# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2727 XNOR2X1_53/a_18_54# XNOR2X1_53/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2728 XNOR2X1_53/a_35_6# XNOR2X1_53/a_2_6# NOR2X1_26/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2729 XNOR2X1_53/a_18_6# XNOR2X1_53/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2730 vdd INVX2_41/Y XNOR2X1_53/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2731 vdd INVX2_31/A XNOR2X1_53/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2732 NOR2X1_26/B XNOR2X1_53/a_2_6# XNOR2X1_53/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2733 XNOR2X1_53/a_35_54# INVX2_41/Y NOR2X1_26/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2734 XNOR2X1_53/a_12_41# INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2735 gnd INVX2_31/A XNOR2X1_53/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2736 gnd INVX2_40/Y XNOR2X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2737 NOR2X1_22/A INVX2_40/Y XNOR2X1_42/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2738 XNOR2X1_42/a_12_41# INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2739 XNOR2X1_42/a_18_54# XNOR2X1_42/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2740 XNOR2X1_42/a_35_6# XNOR2X1_42/a_2_6# NOR2X1_22/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2741 XNOR2X1_42/a_18_6# XNOR2X1_42/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2742 vdd INVX2_40/Y XNOR2X1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2743 vdd INVX2_29/A XNOR2X1_42/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2744 NOR2X1_22/A XNOR2X1_42/a_2_6# XNOR2X1_42/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2745 XNOR2X1_42/a_35_54# INVX2_40/Y NOR2X1_22/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2746 XNOR2X1_42/a_12_41# INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2747 gnd INVX2_29/A XNOR2X1_42/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2748 gnd INVX2_46/A XNOR2X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2749 XNOR2X1_86/Y INVX2_46/A XNOR2X1_86/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2750 XNOR2X1_86/a_12_41# INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2751 XNOR2X1_86/a_18_54# XNOR2X1_86/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2752 XNOR2X1_86/a_35_6# XNOR2X1_86/a_2_6# XNOR2X1_86/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2753 XNOR2X1_86/a_18_6# XNOR2X1_86/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2754 vdd INVX2_46/A XNOR2X1_86/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2755 vdd INVX2_26/A XNOR2X1_86/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2756 XNOR2X1_86/Y XNOR2X1_86/a_2_6# XNOR2X1_86/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2757 XNOR2X1_86/a_35_54# INVX2_46/A XNOR2X1_86/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2758 XNOR2X1_86/a_12_41# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2759 gnd INVX2_26/A XNOR2X1_86/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2760 gnd INVX2_34/A OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2761 vdd DFFSR_7/S INVX2_67/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2762 INVX2_67/A DFFSR_7/S OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2763 INVX2_67/A OAI21X1_4/B OAI21X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2764 OAI21X1_4/a_9_54# INVX2_34/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2765 OAI21X1_4/a_2_6# OAI21X1_4/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2766 DFFNEGX1_2/a_76_6# INVX2_101/Y DFFNEGX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2767 gnd INVX2_101/Y DFFNEGX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2768 DFFNEGX1_2/a_66_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2769 NAND2X1_3/A DFFNEGX1_2/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2770 DFFNEGX1_2/a_23_6# INVX2_101/Y DFFNEGX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2771 DFFNEGX1_2/a_23_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2772 gnd DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2773 vdd DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2774 DFFNEGX1_2/a_61_74# DFFNEGX1_2/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2775 DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2776 DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2777 vdd NAND2X1_3/A DFFNEGX1_2/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2778 gnd NAND2X1_3/A DFFNEGX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2779 DFFNEGX1_2/a_61_6# DFFNEGX1_2/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2780 DFFNEGX1_2/a_76_84# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2781 NAND2X1_3/A DFFNEGX1_2/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2782 vdd INVX2_101/Y DFFNEGX1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2783 DFFNEGX1_2/a_31_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2784 DFFNEGX1_2/a_66_6# INVX2_101/Y DFFNEGX1_2/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2785 DFFNEGX1_2/a_17_74# INVX2_75/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2786 DFFNEGX1_2/a_31_74# INVX2_101/Y DFFNEGX1_2/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2787 DFFNEGX1_2/a_17_6# INVX2_75/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2788 gnd MUX2X1_8/A MUX2X1_8/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2789 MUX2X1_8/a_17_50# INVX2_5/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2790 MUX2X1_8/Y MUX2X1_9/S MUX2X1_8/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2791 MUX2X1_8/a_30_54# MUX2X1_8/a_2_10# MUX2X1_8/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2792 MUX2X1_8/a_17_10# INVX2_5/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2793 vdd MUX2X1_9/S MUX2X1_8/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2794 MUX2X1_8/a_30_10# MUX2X1_9/S MUX2X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2795 gnd MUX2X1_9/S MUX2X1_8/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2796 vdd MUX2X1_8/A MUX2X1_8/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2797 MUX2X1_8/Y MUX2X1_8/a_2_10# MUX2X1_8/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2798 INVX2_61/A NAND3X1_8/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2799 NAND3X1_8/a_9_6# NAND3X1_8/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2800 INVX2_61/A INVX2_43/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2801 INVX2_61/A INVX2_43/Y NAND3X1_8/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2802 vdd NAND3X1_8/B INVX2_61/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2803 NAND3X1_8/a_14_6# NAND3X1_8/B NAND3X1_8/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2804 INVX2_2/Y INVX2_2/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2805 INVX2_2/Y INVX2_2/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2806 AOI21X1_2/a_2_54# AOI21X1_2/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M2807 AOI21X1_2/a_12_6# INVX2_21/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2808 gnd INVX2_66/Y AOI21X1_2/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M2809 vdd INVX2_21/A AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2810 AOI21X1_2/Y INVX2_66/Y AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2811 AOI21X1_2/Y AOI21X1_2/B AOI21X1_2/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2812 gnd NAND2X1_3/A XNOR2X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2813 NAND2X1_9/B NAND2X1_3/A XNOR2X1_10/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2814 XNOR2X1_10/a_12_41# INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2815 XNOR2X1_10/a_18_54# XNOR2X1_10/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2816 XNOR2X1_10/a_35_6# XNOR2X1_10/a_2_6# NAND2X1_9/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2817 XNOR2X1_10/a_18_6# XNOR2X1_10/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2818 vdd NAND2X1_3/A XNOR2X1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2819 vdd INVX2_29/A XNOR2X1_10/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2820 NAND2X1_9/B XNOR2X1_10/a_2_6# XNOR2X1_10/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2821 XNOR2X1_10/a_35_54# NAND2X1_3/A NAND2X1_9/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2822 XNOR2X1_10/a_12_41# INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2823 gnd INVX2_29/A XNOR2X1_10/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2824 gnd NAND2X1_2/A XNOR2X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2825 NAND3X1_5/A NAND2X1_2/A XNOR2X1_21/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2826 XNOR2X1_21/a_12_41# INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2827 XNOR2X1_21/a_18_54# XNOR2X1_21/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2828 XNOR2X1_21/a_35_6# XNOR2X1_21/a_2_6# NAND3X1_5/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2829 XNOR2X1_21/a_18_6# XNOR2X1_21/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2830 vdd NAND2X1_2/A XNOR2X1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2831 vdd INVX2_26/A XNOR2X1_21/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2832 NAND3X1_5/A XNOR2X1_21/a_2_6# XNOR2X1_21/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2833 XNOR2X1_21/a_35_54# NAND2X1_2/A NAND3X1_5/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2834 XNOR2X1_21/a_12_41# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2835 gnd INVX2_26/A XNOR2X1_21/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2836 gnd INVX2_49/Y XNOR2X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2837 NOR2X1_31/A INVX2_49/Y XNOR2X1_76/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2838 XNOR2X1_76/a_12_41# INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2839 XNOR2X1_76/a_18_54# XNOR2X1_76/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2840 XNOR2X1_76/a_35_6# XNOR2X1_76/a_2_6# NOR2X1_31/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2841 XNOR2X1_76/a_18_6# XNOR2X1_76/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2842 vdd INVX2_49/Y XNOR2X1_76/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2843 vdd INVX2_33/A XNOR2X1_76/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2844 NOR2X1_31/A XNOR2X1_76/a_2_6# XNOR2X1_76/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2845 XNOR2X1_76/a_35_54# INVX2_49/Y NOR2X1_31/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2846 XNOR2X1_76/a_12_41# INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2847 gnd INVX2_33/A XNOR2X1_76/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2848 gnd INVX2_45/A XNOR2X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2849 XNOR2X1_43/Y INVX2_45/A XNOR2X1_43/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2850 XNOR2X1_43/a_12_41# INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2851 XNOR2X1_43/a_18_54# XNOR2X1_43/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2852 XNOR2X1_43/a_35_6# XNOR2X1_43/a_2_6# XNOR2X1_43/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2853 XNOR2X1_43/a_18_6# XNOR2X1_43/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2854 vdd INVX2_45/A XNOR2X1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2855 vdd INVX2_29/A XNOR2X1_43/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2856 XNOR2X1_43/Y XNOR2X1_43/a_2_6# XNOR2X1_43/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2857 XNOR2X1_43/a_35_54# INVX2_45/A XNOR2X1_43/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2858 XNOR2X1_43/a_12_41# INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2859 gnd INVX2_29/A XNOR2X1_43/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2860 gnd INVX2_37/A XNOR2X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2861 XNOR2X1_32/Y INVX2_37/A XNOR2X1_32/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2862 XNOR2X1_32/a_12_41# INVX2_46/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2863 XNOR2X1_32/a_18_54# XNOR2X1_32/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2864 XNOR2X1_32/a_35_6# XNOR2X1_32/a_2_6# XNOR2X1_32/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2865 XNOR2X1_32/a_18_6# XNOR2X1_32/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2866 vdd INVX2_37/A XNOR2X1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2867 vdd INVX2_46/A XNOR2X1_32/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2868 XNOR2X1_32/Y XNOR2X1_32/a_2_6# XNOR2X1_32/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2869 XNOR2X1_32/a_35_54# INVX2_37/A XNOR2X1_32/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2870 XNOR2X1_32/a_12_41# INVX2_46/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2871 gnd INVX2_46/A XNOR2X1_32/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2872 gnd INVX2_42/Y XNOR2X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2873 NOR2X1_34/B INVX2_42/Y XNOR2X1_87/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2874 XNOR2X1_87/a_12_41# INVX2_38/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2875 XNOR2X1_87/a_18_54# XNOR2X1_87/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2876 XNOR2X1_87/a_35_6# XNOR2X1_87/a_2_6# NOR2X1_34/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2877 XNOR2X1_87/a_18_6# XNOR2X1_87/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2878 vdd INVX2_42/Y XNOR2X1_87/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2879 vdd INVX2_38/A XNOR2X1_87/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2880 NOR2X1_34/B XNOR2X1_87/a_2_6# XNOR2X1_87/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2881 XNOR2X1_87/a_35_54# INVX2_42/Y NOR2X1_34/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2882 XNOR2X1_87/a_12_41# INVX2_38/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2883 gnd INVX2_38/A XNOR2X1_87/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2884 gnd INVX2_41/Y XNOR2X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2885 NOR2X1_30/B INVX2_41/Y XNOR2X1_65/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2886 XNOR2X1_65/a_12_41# INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2887 XNOR2X1_65/a_18_54# XNOR2X1_65/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2888 XNOR2X1_65/a_35_6# XNOR2X1_65/a_2_6# NOR2X1_30/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2889 XNOR2X1_65/a_18_6# XNOR2X1_65/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2890 vdd INVX2_41/Y XNOR2X1_65/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2891 vdd INVX2_26/A XNOR2X1_65/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2892 NOR2X1_30/B XNOR2X1_65/a_2_6# XNOR2X1_65/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2893 XNOR2X1_65/a_35_54# INVX2_41/Y NOR2X1_30/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2894 XNOR2X1_65/a_12_41# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2895 gnd INVX2_26/A XNOR2X1_65/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2896 gnd INVX2_40/Y XNOR2X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2897 NOR2X1_26/A INVX2_40/Y XNOR2X1_54/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2898 XNOR2X1_54/a_12_41# INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2899 XNOR2X1_54/a_18_54# XNOR2X1_54/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2900 XNOR2X1_54/a_35_6# XNOR2X1_54/a_2_6# NOR2X1_26/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2901 XNOR2X1_54/a_18_6# XNOR2X1_54/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2902 vdd INVX2_40/Y XNOR2X1_54/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2903 vdd INVX2_32/A XNOR2X1_54/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2904 NOR2X1_26/A XNOR2X1_54/a_2_6# XNOR2X1_54/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2905 XNOR2X1_54/a_35_54# INVX2_40/Y NOR2X1_26/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2906 XNOR2X1_54/a_12_41# INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2907 gnd INVX2_32/A XNOR2X1_54/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2908 NOR2X1_0/Y NOR2X1_0/A gnd Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M2909 NOR2X1_0/Y NOR2X1_0/B NOR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M2910 NOR2X1_0/a_9_54# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M2911 gnd NOR2X1_0/B NOR2X1_0/Y Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M2912 gnd OAI21X1_5/A OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2913 vdd DFFSR_7/S INVX2_68/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2914 INVX2_68/A DFFSR_7/S OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2915 INVX2_68/A OAI21X1_5/B OAI21X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2916 OAI21X1_5/a_9_54# OAI21X1_5/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2917 OAI21X1_5/a_2_6# OAI21X1_5/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2918 DFFNEGX1_3/a_76_6# INVX2_101/Y DFFNEGX1_3/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2919 gnd INVX2_101/Y DFFNEGX1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2920 DFFNEGX1_3/a_66_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2921 NAND2X1_4/A DFFNEGX1_3/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2922 DFFNEGX1_3/a_23_6# INVX2_101/Y DFFNEGX1_3/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2923 DFFNEGX1_3/a_23_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2924 gnd DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2925 vdd DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2926 DFFNEGX1_3/a_61_74# DFFNEGX1_3/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2927 DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2928 DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2929 vdd NAND2X1_4/A DFFNEGX1_3/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2930 gnd NAND2X1_4/A DFFNEGX1_3/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2931 DFFNEGX1_3/a_61_6# DFFNEGX1_3/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2932 DFFNEGX1_3/a_76_84# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2933 NAND2X1_4/A DFFNEGX1_3/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2934 vdd INVX2_101/Y DFFNEGX1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2935 DFFNEGX1_3/a_31_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2936 DFFNEGX1_3/a_66_6# INVX2_101/Y DFFNEGX1_3/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2937 DFFNEGX1_3/a_17_74# INVX2_74/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2938 DFFNEGX1_3/a_31_74# INVX2_101/Y DFFNEGX1_3/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2939 DFFNEGX1_3/a_17_6# INVX2_74/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2940 gnd MUX2X1_9/A MUX2X1_9/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2941 MUX2X1_9/a_17_50# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2942 INVX2_8/A MUX2X1_9/S MUX2X1_9/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2943 MUX2X1_9/a_30_54# MUX2X1_9/a_2_10# INVX2_8/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2944 MUX2X1_9/a_17_10# INVX2_6/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2945 vdd MUX2X1_9/S MUX2X1_9/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2946 MUX2X1_9/a_30_10# MUX2X1_9/S INVX2_8/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2947 gnd MUX2X1_9/S MUX2X1_9/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2948 vdd MUX2X1_9/A MUX2X1_9/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2949 INVX2_8/A MUX2X1_9/a_2_10# MUX2X1_9/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2950 INVX2_53/A NAND3X1_9/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M2951 NAND3X1_9/a_9_6# NAND3X1_9/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M2952 INVX2_53/A NOR2X1_31/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2953 INVX2_53/A NOR2X1_31/Y NAND3X1_9/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M2954 vdd NAND3X1_9/B INVX2_53/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2955 NAND3X1_9/a_14_6# NAND3X1_9/B NAND3X1_9/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M2956 INVX2_3/Y INVX2_3/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2957 INVX2_3/Y INVX2_3/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2958 AOI21X1_3/a_2_54# AOI21X1_3/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M2959 AOI21X1_3/a_12_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2960 gnd NOR2X1_35/Y INVX2_64/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M2961 vdd NOR2X1_36/Y AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2962 INVX2_64/A NOR2X1_35/Y AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2963 INVX2_64/A AOI21X1_3/B AOI21X1_3/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2964 gnd NAND2X1_2/A XNOR2X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2965 NAND2X1_9/A NAND2X1_2/A XNOR2X1_11/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2966 XNOR2X1_11/a_12_41# INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2967 XNOR2X1_11/a_18_54# XNOR2X1_11/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2968 XNOR2X1_11/a_35_6# XNOR2X1_11/a_2_6# NAND2X1_9/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2969 XNOR2X1_11/a_18_6# XNOR2X1_11/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2970 vdd NAND2X1_2/A XNOR2X1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2971 vdd INVX2_28/A XNOR2X1_11/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2972 NAND2X1_9/A XNOR2X1_11/a_2_6# XNOR2X1_11/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2973 XNOR2X1_11/a_35_54# NAND2X1_2/A NAND2X1_9/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2974 XNOR2X1_11/a_12_41# INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2975 gnd INVX2_28/A XNOR2X1_11/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2976 gnd INVX2_45/A XNOR2X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2977 XNOR2X1_55/Y INVX2_45/A XNOR2X1_55/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2978 XNOR2X1_55/a_12_41# INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2979 XNOR2X1_55/a_18_54# XNOR2X1_55/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2980 XNOR2X1_55/a_35_6# XNOR2X1_55/a_2_6# XNOR2X1_55/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2981 XNOR2X1_55/a_18_6# XNOR2X1_55/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2982 vdd INVX2_45/A XNOR2X1_55/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2983 vdd INVX2_32/A XNOR2X1_55/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2984 XNOR2X1_55/Y XNOR2X1_55/a_2_6# XNOR2X1_55/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2985 XNOR2X1_55/a_35_54# INVX2_45/A XNOR2X1_55/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2986 XNOR2X1_55/a_12_41# INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2987 gnd INVX2_32/A XNOR2X1_55/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2988 gnd XNOR2X1_22/A XNOR2X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2989 out_Bnum[1] XNOR2X1_22/A XNOR2X1_22/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2990 XNOR2X1_22/a_12_41# INVX2_58/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2991 XNOR2X1_22/a_18_54# XNOR2X1_22/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2992 XNOR2X1_22/a_35_6# XNOR2X1_22/a_2_6# out_Bnum[1] Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2993 XNOR2X1_22/a_18_6# XNOR2X1_22/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2994 vdd XNOR2X1_22/A XNOR2X1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2995 vdd INVX2_58/Y XNOR2X1_22/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2996 out_Bnum[1] XNOR2X1_22/a_2_6# XNOR2X1_22/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2997 XNOR2X1_22/a_35_54# XNOR2X1_22/A out_Bnum[1] vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2998 XNOR2X1_22/a_12_41# INVX2_58/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2999 gnd INVX2_58/Y XNOR2X1_22/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3000 gnd INVX2_35/A XNOR2X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3001 XNOR2X1_33/Y INVX2_35/A XNOR2X1_33/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3002 XNOR2X1_33/a_12_41# INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3003 XNOR2X1_33/a_18_54# XNOR2X1_33/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3004 XNOR2X1_33/a_35_6# XNOR2X1_33/a_2_6# XNOR2X1_33/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3005 XNOR2X1_33/a_18_6# XNOR2X1_33/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3006 vdd INVX2_35/A XNOR2X1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3007 vdd INVX2_44/A XNOR2X1_33/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3008 XNOR2X1_33/Y XNOR2X1_33/a_2_6# XNOR2X1_33/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3009 XNOR2X1_33/a_35_54# INVX2_35/A XNOR2X1_33/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3010 XNOR2X1_33/a_12_41# INVX2_44/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3011 gnd INVX2_44/A XNOR2X1_33/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3012 gnd INVX2_50/A XNOR2X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3013 NAND3X1_9/B INVX2_50/A XNOR2X1_77/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3014 XNOR2X1_77/a_12_41# INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3015 XNOR2X1_77/a_18_54# XNOR2X1_77/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3016 XNOR2X1_77/a_35_6# XNOR2X1_77/a_2_6# NAND3X1_9/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3017 XNOR2X1_77/a_18_6# XNOR2X1_77/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3018 vdd INVX2_50/A XNOR2X1_77/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3019 vdd INVX2_32/A XNOR2X1_77/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3020 NAND3X1_9/B XNOR2X1_77/a_2_6# XNOR2X1_77/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3021 XNOR2X1_77/a_35_54# INVX2_50/A NAND3X1_9/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3022 XNOR2X1_77/a_12_41# INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3023 gnd INVX2_32/A XNOR2X1_77/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3024 gnd INVX2_46/A XNOR2X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3025 XNOR2X1_44/Y INVX2_46/A XNOR2X1_44/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3026 XNOR2X1_44/a_12_41# INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3027 XNOR2X1_44/a_18_54# XNOR2X1_44/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3028 XNOR2X1_44/a_35_6# XNOR2X1_44/a_2_6# XNOR2X1_44/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3029 XNOR2X1_44/a_18_6# XNOR2X1_44/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3030 vdd INVX2_46/A XNOR2X1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3031 vdd INVX2_28/A XNOR2X1_44/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3032 XNOR2X1_44/Y XNOR2X1_44/a_2_6# XNOR2X1_44/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3033 XNOR2X1_44/a_35_54# INVX2_46/A XNOR2X1_44/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3034 XNOR2X1_44/a_12_41# INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3035 gnd INVX2_28/A XNOR2X1_44/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3036 gnd INVX2_39/Y XNOR2X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3037 NOR2X1_34/A INVX2_39/Y XNOR2X1_88/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3038 XNOR2X1_88/a_12_41# INVX2_35/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3039 XNOR2X1_88/a_18_54# XNOR2X1_88/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3040 XNOR2X1_88/a_35_6# XNOR2X1_88/a_2_6# NOR2X1_34/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3041 XNOR2X1_88/a_18_6# XNOR2X1_88/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3042 vdd INVX2_39/Y XNOR2X1_88/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3043 vdd INVX2_35/A XNOR2X1_88/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3044 NOR2X1_34/A XNOR2X1_88/a_2_6# XNOR2X1_88/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3045 XNOR2X1_88/a_35_54# INVX2_39/Y NOR2X1_34/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3046 XNOR2X1_88/a_12_41# INVX2_35/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3047 gnd INVX2_35/A XNOR2X1_88/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3048 gnd INVX2_40/Y XNOR2X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3049 NOR2X1_30/A INVX2_40/Y XNOR2X1_66/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3050 XNOR2X1_66/a_12_41# INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3051 XNOR2X1_66/a_18_54# XNOR2X1_66/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3052 XNOR2X1_66/a_35_6# XNOR2X1_66/a_2_6# NOR2X1_30/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3053 XNOR2X1_66/a_18_6# XNOR2X1_66/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3054 vdd INVX2_40/Y XNOR2X1_66/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3055 vdd INVX2_25/A XNOR2X1_66/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3056 NOR2X1_30/A XNOR2X1_66/a_2_6# XNOR2X1_66/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3057 XNOR2X1_66/a_35_54# INVX2_40/Y NOR2X1_30/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3058 XNOR2X1_66/a_12_41# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3059 gnd INVX2_25/A XNOR2X1_66/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3060 NOR2X1_1/Y INVX2_9/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3061 NOR2X1_1/Y NOR2X1_1/B NOR2X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3062 NOR2X1_1/a_9_54# INVX2_9/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3063 gnd NOR2X1_1/B NOR2X1_1/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3064 gnd INVX2_70/Y OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3065 vdd DFFSR_7/S INVX2_71/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3066 INVX2_71/A DFFSR_7/S OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3067 INVX2_71/A OAI21X1_6/B OAI21X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3068 OAI21X1_6/a_9_54# INVX2_70/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3069 OAI21X1_6/a_2_6# OAI21X1_6/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3070 gnd OAI22X1_6/A OAI22X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3071 OAI22X1_30/a_2_6# INVX2_98/Y OAI22X1_30/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3072 OAI22X1_30/Y INVX2_89/Y OAI22X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3073 OAI22X1_30/Y INVX2_49/Y OAI22X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3074 OAI22X1_30/a_28_54# INVX2_89/Y OAI22X1_30/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3075 OAI22X1_30/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3076 OAI22X1_30/a_2_6# INVX2_49/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3077 vdd INVX2_98/Y OAI22X1_30/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3078 DFFNEGX1_4/a_76_6# INVX2_101/Y DFFNEGX1_4/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3079 gnd INVX2_101/Y DFFNEGX1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3080 DFFNEGX1_4/a_66_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3081 INVX2_18/A DFFNEGX1_4/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3082 DFFNEGX1_4/a_23_6# INVX2_101/Y DFFNEGX1_4/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3083 DFFNEGX1_4/a_23_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3084 gnd DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3085 vdd DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3086 DFFNEGX1_4/a_61_74# DFFNEGX1_4/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3087 DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3088 DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3089 vdd INVX2_18/A DFFNEGX1_4/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3090 gnd INVX2_18/A DFFNEGX1_4/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3091 DFFNEGX1_4/a_61_6# DFFNEGX1_4/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3092 DFFNEGX1_4/a_76_84# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3093 INVX2_18/A DFFNEGX1_4/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3094 vdd INVX2_101/Y DFFNEGX1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3095 DFFNEGX1_4/a_31_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3096 DFFNEGX1_4/a_66_6# INVX2_101/Y DFFNEGX1_4/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3097 DFFNEGX1_4/a_17_74# OAI22X1_22/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3098 DFFNEGX1_4/a_31_74# INVX2_101/Y DFFNEGX1_4/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3099 DFFNEGX1_4/a_17_6# OAI22X1_22/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3100 INVX2_4/Y INVX2_4/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3101 INVX2_4/Y INVX2_4/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3102 gnd NAND2X1_4/A XNOR2X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3103 XNOR2X1_12/Y NAND2X1_4/A XNOR2X1_12/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3104 XNOR2X1_12/a_12_41# INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3105 XNOR2X1_12/a_18_54# XNOR2X1_12/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3106 XNOR2X1_12/a_35_6# XNOR2X1_12/a_2_6# XNOR2X1_12/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3107 XNOR2X1_12/a_18_6# XNOR2X1_12/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3108 vdd NAND2X1_4/A XNOR2X1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3109 vdd INVX2_30/A XNOR2X1_12/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3110 XNOR2X1_12/Y XNOR2X1_12/a_2_6# XNOR2X1_12/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3111 XNOR2X1_12/a_35_54# NAND2X1_4/A XNOR2X1_12/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3112 XNOR2X1_12/a_12_41# INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3113 gnd INVX2_30/A XNOR2X1_12/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3114 gnd INVX2_52/Y XNOR2X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3115 NOR2X1_15/B INVX2_52/Y XNOR2X1_23/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3116 XNOR2X1_23/a_12_41# INVX2_38/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3117 XNOR2X1_23/a_18_54# XNOR2X1_23/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3118 XNOR2X1_23/a_35_6# XNOR2X1_23/a_2_6# NOR2X1_15/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3119 XNOR2X1_23/a_18_6# XNOR2X1_23/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3120 vdd INVX2_52/Y XNOR2X1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3121 vdd INVX2_38/A XNOR2X1_23/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3122 NOR2X1_15/B XNOR2X1_23/a_2_6# XNOR2X1_23/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3123 XNOR2X1_23/a_35_54# INVX2_52/Y NOR2X1_15/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3124 XNOR2X1_23/a_12_41# INVX2_38/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3125 gnd INVX2_38/A XNOR2X1_23/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3126 gnd INVX2_46/A XNOR2X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3127 XNOR2X1_56/Y INVX2_46/A XNOR2X1_56/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3128 XNOR2X1_56/a_12_41# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3129 XNOR2X1_56/a_18_54# XNOR2X1_56/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3130 XNOR2X1_56/a_35_6# XNOR2X1_56/a_2_6# XNOR2X1_56/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3131 XNOR2X1_56/a_18_6# XNOR2X1_56/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3132 vdd INVX2_46/A XNOR2X1_56/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3133 vdd INVX2_31/A XNOR2X1_56/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3134 XNOR2X1_56/Y XNOR2X1_56/a_2_6# XNOR2X1_56/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3135 XNOR2X1_56/a_35_54# INVX2_46/A XNOR2X1_56/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3136 XNOR2X1_56/a_12_41# INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3137 gnd INVX2_31/A XNOR2X1_56/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3138 gnd INVX2_38/A XNOR2X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3139 XNOR2X1_34/Y INVX2_38/A XNOR2X1_34/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3140 XNOR2X1_34/a_12_41# INVX2_47/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3141 XNOR2X1_34/a_18_54# XNOR2X1_34/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3142 XNOR2X1_34/a_35_6# XNOR2X1_34/a_2_6# XNOR2X1_34/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3143 XNOR2X1_34/a_18_6# XNOR2X1_34/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3144 vdd INVX2_38/A XNOR2X1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3145 vdd INVX2_47/A XNOR2X1_34/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3146 XNOR2X1_34/Y XNOR2X1_34/a_2_6# XNOR2X1_34/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3147 XNOR2X1_34/a_35_54# INVX2_38/A XNOR2X1_34/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3148 XNOR2X1_34/a_12_41# INVX2_47/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3149 gnd INVX2_47/A XNOR2X1_34/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3150 gnd INVX2_44/A XNOR2X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3151 XNOR2X1_45/Y INVX2_44/A XNOR2X1_45/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3152 XNOR2X1_45/a_12_41# INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3153 XNOR2X1_45/a_18_54# XNOR2X1_45/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3154 XNOR2X1_45/a_35_6# XNOR2X1_45/a_2_6# XNOR2X1_45/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3155 XNOR2X1_45/a_18_6# XNOR2X1_45/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3156 vdd INVX2_44/A XNOR2X1_45/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3157 vdd INVX2_30/A XNOR2X1_45/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3158 XNOR2X1_45/Y XNOR2X1_45/a_2_6# XNOR2X1_45/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3159 XNOR2X1_45/a_35_54# INVX2_44/A XNOR2X1_45/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3160 XNOR2X1_45/a_12_41# INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3161 gnd INVX2_30/A XNOR2X1_45/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3162 gnd INVX2_50/A XNOR2X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3163 XNOR2X1_67/Y INVX2_50/A XNOR2X1_67/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3164 XNOR2X1_67/a_12_41# INVX2_25/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3165 XNOR2X1_67/a_18_54# XNOR2X1_67/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3166 XNOR2X1_67/a_35_6# XNOR2X1_67/a_2_6# XNOR2X1_67/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3167 XNOR2X1_67/a_18_6# XNOR2X1_67/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3168 vdd INVX2_50/A XNOR2X1_67/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3169 vdd INVX2_25/A XNOR2X1_67/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3170 XNOR2X1_67/Y XNOR2X1_67/a_2_6# XNOR2X1_67/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3171 XNOR2X1_67/a_35_54# INVX2_50/A XNOR2X1_67/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3172 XNOR2X1_67/a_12_41# INVX2_25/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3173 gnd INVX2_25/A XNOR2X1_67/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3174 gnd INVX2_51/A XNOR2X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3175 NAND3X1_9/A INVX2_51/A XNOR2X1_78/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3176 XNOR2X1_78/a_12_41# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3177 XNOR2X1_78/a_18_54# XNOR2X1_78/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3178 XNOR2X1_78/a_35_6# XNOR2X1_78/a_2_6# NAND3X1_9/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3179 XNOR2X1_78/a_18_6# XNOR2X1_78/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3180 vdd INVX2_51/A XNOR2X1_78/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3181 vdd INVX2_31/A XNOR2X1_78/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3182 NAND3X1_9/A XNOR2X1_78/a_2_6# XNOR2X1_78/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3183 XNOR2X1_78/a_35_54# INVX2_51/A NAND3X1_9/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3184 XNOR2X1_78/a_12_41# INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3185 gnd INVX2_31/A XNOR2X1_78/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3186 gnd INVX2_36/A XNOR2X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3187 XNOR2X1_89/Y INVX2_36/A XNOR2X1_89/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3188 XNOR2X1_89/a_12_41# INVX2_40/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3189 XNOR2X1_89/a_18_54# XNOR2X1_89/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3190 XNOR2X1_89/a_35_6# XNOR2X1_89/a_2_6# XNOR2X1_89/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3191 XNOR2X1_89/a_18_6# XNOR2X1_89/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3192 vdd INVX2_36/A XNOR2X1_89/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3193 vdd INVX2_40/A XNOR2X1_89/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3194 XNOR2X1_89/Y XNOR2X1_89/a_2_6# XNOR2X1_89/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3195 XNOR2X1_89/a_35_54# INVX2_36/A XNOR2X1_89/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3196 XNOR2X1_89/a_12_41# INVX2_40/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3197 gnd INVX2_40/A XNOR2X1_89/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3198 NOR2X1_2/Y INVX2_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3199 NOR2X1_2/Y INVX2_7/Y NOR2X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3200 NOR2X1_2/a_9_54# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3201 gnd INVX2_7/Y NOR2X1_2/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3202 gnd INVX2_70/Y OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3203 vdd OAI21X1_7/C OAI21X1_7/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3204 OAI21X1_7/Y OAI21X1_7/C OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3205 OAI21X1_7/Y OAI21X1_7/B OAI21X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3206 OAI21X1_7/a_9_54# INVX2_70/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3207 OAI21X1_7/a_2_6# OAI21X1_7/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3208 gnd INVX2_24/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3209 OAI22X1_20/a_2_6# INVX2_71/Y OAI22X1_20/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3210 OAI22X1_20/Y NAND2X1_4/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3211 OAI22X1_20/Y INVX2_71/A OAI22X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3212 OAI22X1_20/a_28_54# NAND2X1_4/Y OAI22X1_20/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3213 OAI22X1_20/a_9_54# INVX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3214 OAI22X1_20/a_2_6# INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3215 vdd INVX2_71/Y OAI22X1_20/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3216 gnd OAI22X1_6/A OAI22X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3217 OAI22X1_31/a_2_6# INVX2_98/Y OAI22X1_31/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3218 OAI22X1_31/Y INVX2_90/Y OAI22X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3219 OAI22X1_31/Y INVX2_47/Y OAI22X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3220 OAI22X1_31/a_28_54# INVX2_90/Y OAI22X1_31/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3221 OAI22X1_31/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3222 OAI22X1_31/a_2_6# INVX2_47/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3223 vdd INVX2_98/Y OAI22X1_31/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3224 DFFNEGX1_5/a_76_6# INVX2_101/Y DFFNEGX1_5/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3225 gnd INVX2_101/Y DFFNEGX1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3226 DFFNEGX1_5/a_66_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3227 INVX2_19/A DFFNEGX1_5/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3228 DFFNEGX1_5/a_23_6# INVX2_101/Y DFFNEGX1_5/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3229 DFFNEGX1_5/a_23_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3230 gnd DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3231 vdd DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3232 DFFNEGX1_5/a_61_74# DFFNEGX1_5/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3233 DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3234 DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3235 vdd INVX2_19/A DFFNEGX1_5/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3236 gnd INVX2_19/A DFFNEGX1_5/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3237 DFFNEGX1_5/a_61_6# DFFNEGX1_5/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3238 DFFNEGX1_5/a_76_84# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3239 INVX2_19/A DFFNEGX1_5/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3240 vdd INVX2_101/Y DFFNEGX1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3241 DFFNEGX1_5/a_31_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3242 DFFNEGX1_5/a_66_6# INVX2_101/Y DFFNEGX1_5/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3243 DFFNEGX1_5/a_17_74# OAI21X1_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3244 DFFNEGX1_5/a_31_74# INVX2_101/Y DFFNEGX1_5/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3245 DFFNEGX1_5/a_17_6# OAI21X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3246 OAI21X1_4/B INVX2_70/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3247 NAND2X1_0/a_9_6# INVX2_70/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3248 vdd NOR2X1_8/Y OAI21X1_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3249 OAI21X1_4/B NOR2X1_8/Y NAND2X1_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3250 INVX2_5/Y INVX2_5/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3251 INVX2_5/Y INVX2_5/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3252 gnd AOI22X1_3/C XNOR2X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3253 XNOR2X1_13/Y AOI22X1_3/C XNOR2X1_13/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3254 XNOR2X1_13/a_12_41# INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3255 XNOR2X1_13/a_18_54# XNOR2X1_13/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3256 XNOR2X1_13/a_35_6# XNOR2X1_13/a_2_6# XNOR2X1_13/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3257 XNOR2X1_13/a_18_6# XNOR2X1_13/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3258 vdd AOI22X1_3/C XNOR2X1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3259 vdd INVX2_27/A XNOR2X1_13/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3260 XNOR2X1_13/Y XNOR2X1_13/a_2_6# XNOR2X1_13/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3261 XNOR2X1_13/a_35_54# AOI22X1_3/C XNOR2X1_13/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3262 XNOR2X1_13/a_12_41# INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3263 gnd INVX2_27/A XNOR2X1_13/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3264 gnd INVX2_44/A XNOR2X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3265 XNOR2X1_57/Y INVX2_44/A XNOR2X1_57/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3266 XNOR2X1_57/a_12_41# INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3267 XNOR2X1_57/a_18_54# XNOR2X1_57/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3268 XNOR2X1_57/a_35_6# XNOR2X1_57/a_2_6# XNOR2X1_57/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3269 XNOR2X1_57/a_18_6# XNOR2X1_57/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3270 vdd INVX2_44/A XNOR2X1_57/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3271 vdd INVX2_33/A XNOR2X1_57/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3272 XNOR2X1_57/Y XNOR2X1_57/a_2_6# XNOR2X1_57/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3273 XNOR2X1_57/a_35_54# INVX2_44/A XNOR2X1_57/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3274 XNOR2X1_57/a_12_41# INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3275 gnd INVX2_33/A XNOR2X1_57/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3276 gnd INVX2_47/A XNOR2X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3277 XNOR2X1_46/Y INVX2_47/A XNOR2X1_46/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3278 XNOR2X1_46/a_12_41# INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3279 XNOR2X1_46/a_18_54# XNOR2X1_46/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3280 XNOR2X1_46/a_35_6# XNOR2X1_46/a_2_6# XNOR2X1_46/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3281 XNOR2X1_46/a_18_6# XNOR2X1_46/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3282 vdd INVX2_47/A XNOR2X1_46/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3283 vdd INVX2_27/A XNOR2X1_46/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3284 XNOR2X1_46/Y XNOR2X1_46/a_2_6# XNOR2X1_46/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3285 XNOR2X1_46/a_35_54# INVX2_47/A XNOR2X1_46/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3286 XNOR2X1_46/a_12_41# INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3287 gnd INVX2_27/A XNOR2X1_46/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3288 gnd INVX2_49/Y XNOR2X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3289 NOR2X1_15/A INVX2_49/Y XNOR2X1_24/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3290 XNOR2X1_24/a_12_41# INVX2_35/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3291 XNOR2X1_24/a_18_54# XNOR2X1_24/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3292 XNOR2X1_24/a_35_6# XNOR2X1_24/a_2_6# NOR2X1_15/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3293 XNOR2X1_24/a_18_6# XNOR2X1_24/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3294 vdd INVX2_49/Y XNOR2X1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3295 vdd INVX2_35/A XNOR2X1_24/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3296 NOR2X1_15/A XNOR2X1_24/a_2_6# XNOR2X1_24/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3297 XNOR2X1_24/a_35_54# INVX2_49/Y NOR2X1_15/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3298 XNOR2X1_24/a_12_41# INVX2_35/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3299 gnd INVX2_35/A XNOR2X1_24/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3300 gnd INVX2_52/Y XNOR2X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3301 NOR2X1_19/B INVX2_52/Y XNOR2X1_35/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3302 XNOR2X1_35/a_12_41# INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3303 XNOR2X1_35/a_18_54# XNOR2X1_35/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3304 XNOR2X1_35/a_35_6# XNOR2X1_35/a_2_6# NOR2X1_19/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3305 XNOR2X1_35/a_18_6# XNOR2X1_35/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3306 vdd INVX2_52/Y XNOR2X1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3307 vdd INVX2_27/A XNOR2X1_35/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3308 NOR2X1_19/B XNOR2X1_35/a_2_6# XNOR2X1_35/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3309 XNOR2X1_35/a_35_54# INVX2_52/Y NOR2X1_19/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3310 XNOR2X1_35/a_12_41# INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3311 gnd INVX2_27/A XNOR2X1_35/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3312 gnd INVX2_51/A XNOR2X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3313 XNOR2X1_68/Y INVX2_51/A XNOR2X1_68/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3314 XNOR2X1_68/a_12_41# INVX2_26/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3315 XNOR2X1_68/a_18_54# XNOR2X1_68/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3316 XNOR2X1_68/a_35_6# XNOR2X1_68/a_2_6# XNOR2X1_68/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3317 XNOR2X1_68/a_18_6# XNOR2X1_68/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3318 vdd INVX2_51/A XNOR2X1_68/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3319 vdd INVX2_26/A XNOR2X1_68/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3320 XNOR2X1_68/Y XNOR2X1_68/a_2_6# XNOR2X1_68/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3321 XNOR2X1_68/a_35_54# INVX2_51/A XNOR2X1_68/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3322 XNOR2X1_68/a_12_41# INVX2_26/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3323 gnd INVX2_26/A XNOR2X1_68/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3324 gnd INVX2_57/Y XNOR2X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3325 NOR2X1_32/B INVX2_57/Y XNOR2X1_79/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3326 XNOR2X1_79/a_12_41# INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3327 XNOR2X1_79/a_18_54# XNOR2X1_79/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3328 XNOR2X1_79/a_35_6# XNOR2X1_79/a_2_6# NOR2X1_32/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3329 XNOR2X1_79/a_18_6# XNOR2X1_79/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3330 vdd INVX2_57/Y XNOR2X1_79/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3331 vdd INVX2_27/A XNOR2X1_79/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3332 NOR2X1_32/B XNOR2X1_79/a_2_6# XNOR2X1_79/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3333 XNOR2X1_79/a_35_54# INVX2_57/Y NOR2X1_32/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3334 XNOR2X1_79/a_12_41# INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3335 gnd INVX2_27/A XNOR2X1_79/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3336 NOR2X1_3/Y INVX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3337 NOR2X1_3/Y INVX2_4/Y NOR2X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3338 NOR2X1_3/a_9_54# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3339 gnd INVX2_4/Y NOR2X1_3/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3340 OR2X1_0/a_2_54# OR2X1_0/A gnd Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M3341 OR2X1_0/Y OR2X1_0/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0.11n ps=46u
M3342 OR2X1_0/Y OR2X1_0/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M3343 vdd OR2X1_0/B OR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=59.999996p ps=43u
M3344 OR2X1_0/a_9_54# OR2X1_0/A OR2X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M3345 gnd OR2X1_0/B OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=29.999998p ps=16u
M3346 gnd NOR2X1_6/A OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3347 vdd OAI21X1_8/C OAI21X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3348 OAI21X1_8/Y OAI21X1_8/C OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3349 OAI21X1_8/Y NOR2X1_8/B OAI21X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3350 OAI21X1_8/a_9_54# NOR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3351 OAI21X1_8/a_2_6# NOR2X1_8/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3352 gnd INVX2_23/Y OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3353 OAI22X1_21/a_2_6# INVX2_71/Y OAI22X1_21/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3354 OAI22X1_21/Y OAI22X1_7/D OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3355 OAI22X1_21/Y INVX2_71/A OAI22X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3356 OAI22X1_21/a_28_54# OAI22X1_7/D OAI22X1_21/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3357 OAI22X1_21/a_9_54# INVX2_23/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3358 OAI22X1_21/a_2_6# INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3359 vdd INVX2_71/Y OAI22X1_21/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3360 gnd INVX2_67/A OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3361 OAI22X1_10/a_2_6# INVX2_67/Y OAI22X1_10/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3362 OAI22X1_10/Y NAND2X1_4/Y OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3363 OAI22X1_10/Y INVX2_35/Y OAI22X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3364 OAI22X1_10/a_28_54# NAND2X1_4/Y OAI22X1_10/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3365 OAI22X1_10/a_9_54# INVX2_67/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3366 OAI22X1_10/a_2_6# INVX2_35/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3367 vdd INVX2_67/Y OAI22X1_10/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3368 gnd XNOR2X1_74/Y OAI22X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3369 OAI22X1_32/a_2_6# INVX2_60/A NAND3X1_8/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3370 NAND3X1_8/B INVX2_53/A OAI22X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3371 NAND3X1_8/B INVX2_48/A OAI22X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3372 OAI22X1_32/a_28_54# INVX2_53/A NAND3X1_8/B vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3373 OAI22X1_32/a_9_54# XNOR2X1_74/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3374 OAI22X1_32/a_2_6# INVX2_48/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3375 vdd INVX2_60/A OAI22X1_32/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3376 DFFNEGX1_6/a_76_6# INVX2_101/Y DFFNEGX1_6/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3377 gnd INVX2_101/Y DFFNEGX1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3378 DFFNEGX1_6/a_66_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3379 OR2X1_0/B DFFNEGX1_6/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3380 DFFNEGX1_6/a_23_6# INVX2_101/Y DFFNEGX1_6/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3381 DFFNEGX1_6/a_23_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3382 gnd DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3383 vdd DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3384 DFFNEGX1_6/a_61_74# DFFNEGX1_6/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3385 DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3386 DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3387 vdd OR2X1_0/B DFFNEGX1_6/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3388 gnd OR2X1_0/B DFFNEGX1_6/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3389 DFFNEGX1_6/a_61_6# DFFNEGX1_6/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3390 DFFNEGX1_6/a_76_84# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3391 OR2X1_0/B DFFNEGX1_6/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3392 vdd INVX2_101/Y DFFNEGX1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3393 DFFNEGX1_6/a_31_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3394 DFFNEGX1_6/a_66_6# INVX2_101/Y DFFNEGX1_6/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3395 DFFNEGX1_6/a_17_74# NOR2X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3396 DFFNEGX1_6/a_31_74# INVX2_101/Y DFFNEGX1_6/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3397 DFFNEGX1_6/a_17_6# NOR2X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3398 OAI21X1_5/B INVX2_19/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3399 NAND2X1_1/a_9_6# INVX2_19/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3400 vdd AND2X2_2/B OAI21X1_5/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3401 OAI21X1_5/B AND2X2_2/B NAND2X1_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3402 INVX2_6/Y INVX2_6/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3403 INVX2_6/Y INVX2_6/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3404 gnd AOI22X1_3/C XNOR2X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3405 NOR2X1_10/B AOI22X1_3/C XNOR2X1_14/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3406 XNOR2X1_14/a_12_41# INVX2_18/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3407 XNOR2X1_14/a_18_54# XNOR2X1_14/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3408 XNOR2X1_14/a_35_6# XNOR2X1_14/a_2_6# NOR2X1_10/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3409 XNOR2X1_14/a_18_6# XNOR2X1_14/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3410 vdd AOI22X1_3/C XNOR2X1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3411 vdd INVX2_18/Y XNOR2X1_14/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3412 NOR2X1_10/B XNOR2X1_14/a_2_6# XNOR2X1_14/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3413 XNOR2X1_14/a_35_54# AOI22X1_3/C NOR2X1_10/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3414 XNOR2X1_14/a_12_41# INVX2_18/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3415 gnd INVX2_18/Y XNOR2X1_14/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3416 gnd INVX2_47/A XNOR2X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3417 XNOR2X1_58/Y INVX2_47/A XNOR2X1_58/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3418 XNOR2X1_58/a_12_41# INVX2_18/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3419 XNOR2X1_58/a_18_54# XNOR2X1_58/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3420 XNOR2X1_58/a_35_6# XNOR2X1_58/a_2_6# XNOR2X1_58/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3421 XNOR2X1_58/a_18_6# XNOR2X1_58/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3422 vdd INVX2_47/A XNOR2X1_58/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3423 vdd INVX2_18/A XNOR2X1_58/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3424 XNOR2X1_58/Y XNOR2X1_58/a_2_6# XNOR2X1_58/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3425 XNOR2X1_58/a_35_54# INVX2_47/A XNOR2X1_58/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3426 XNOR2X1_58/a_12_41# INVX2_18/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3427 gnd INVX2_18/A XNOR2X1_58/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3428 gnd INVX2_49/A XNOR2X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3429 XNOR2X1_69/Y INVX2_49/A XNOR2X1_69/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3430 XNOR2X1_69/a_12_41# INVX2_24/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3431 XNOR2X1_69/a_18_54# XNOR2X1_69/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3432 XNOR2X1_69/a_35_6# XNOR2X1_69/a_2_6# XNOR2X1_69/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3433 XNOR2X1_69/a_18_6# XNOR2X1_69/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3434 vdd INVX2_49/A XNOR2X1_69/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3435 vdd INVX2_24/A XNOR2X1_69/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3436 XNOR2X1_69/Y XNOR2X1_69/a_2_6# XNOR2X1_69/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3437 XNOR2X1_69/a_35_54# INVX2_49/A XNOR2X1_69/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3438 XNOR2X1_69/a_12_41# INVX2_24/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3439 gnd INVX2_24/A XNOR2X1_69/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3440 gnd INVX2_49/Y XNOR2X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3441 NOR2X1_19/A INVX2_49/Y XNOR2X1_36/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3442 XNOR2X1_36/a_12_41# INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3443 XNOR2X1_36/a_18_54# XNOR2X1_36/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3444 XNOR2X1_36/a_35_6# XNOR2X1_36/a_2_6# NOR2X1_19/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3445 XNOR2X1_36/a_18_6# XNOR2X1_36/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3446 vdd INVX2_49/Y XNOR2X1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3447 vdd INVX2_30/A XNOR2X1_36/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3448 NOR2X1_19/A XNOR2X1_36/a_2_6# XNOR2X1_36/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3449 XNOR2X1_36/a_35_54# INVX2_49/Y NOR2X1_19/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3450 XNOR2X1_36/a_12_41# INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3451 gnd INVX2_30/A XNOR2X1_36/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3452 gnd INVX2_51/Y XNOR2X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3453 NOR2X1_16/B INVX2_51/Y XNOR2X1_25/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3454 XNOR2X1_25/a_12_41# INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3455 XNOR2X1_25/a_18_54# XNOR2X1_25/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3456 XNOR2X1_25/a_35_6# XNOR2X1_25/a_2_6# NOR2X1_16/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3457 XNOR2X1_25/a_18_6# XNOR2X1_25/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3458 vdd INVX2_51/Y XNOR2X1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3459 vdd INVX2_37/A XNOR2X1_25/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3460 NOR2X1_16/B XNOR2X1_25/a_2_6# XNOR2X1_25/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3461 XNOR2X1_25/a_35_54# INVX2_51/Y NOR2X1_16/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3462 XNOR2X1_25/a_12_41# INVX2_37/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3463 gnd INVX2_37/A XNOR2X1_25/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3464 gnd INVX2_57/Y XNOR2X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3465 NOR2X1_23/B INVX2_57/Y XNOR2X1_47/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3466 XNOR2X1_47/a_12_41# INVX2_18/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3467 XNOR2X1_47/a_18_54# XNOR2X1_47/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3468 XNOR2X1_47/a_35_6# XNOR2X1_47/a_2_6# NOR2X1_23/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3469 XNOR2X1_47/a_18_6# XNOR2X1_47/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3470 vdd INVX2_57/Y XNOR2X1_47/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3471 vdd INVX2_18/A XNOR2X1_47/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3472 NOR2X1_23/B XNOR2X1_47/a_2_6# XNOR2X1_47/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3473 XNOR2X1_47/a_35_54# INVX2_57/Y NOR2X1_23/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3474 XNOR2X1_47/a_12_41# INVX2_18/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3475 gnd INVX2_18/A XNOR2X1_47/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3476 NOR2X1_5/A DFFSR_7/D gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3477 NOR2X1_5/A INVX2_0/A NOR2X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3478 NOR2X1_4/a_9_54# DFFSR_7/D vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3479 gnd INVX2_0/A NOR2X1_5/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3480 gnd INVX2_73/Y OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3481 vdd OAI21X1_9/C OAI21X1_9/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3482 OAI21X1_9/Y OAI21X1_9/C OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3483 OAI21X1_9/Y NOR2X1_7/A OAI21X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3484 OAI21X1_9/a_9_54# INVX2_73/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3485 OAI21X1_9/a_2_6# NOR2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3486 gnd INVX2_30/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3487 OAI22X1_11/a_2_6# INVX2_68/Y OAI22X1_11/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3488 OAI22X1_11/Y NAND2X1_4/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3489 OAI22X1_11/Y INVX2_68/A OAI22X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3490 OAI22X1_11/a_28_54# NAND2X1_4/Y OAI22X1_11/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3491 OAI22X1_11/a_9_54# INVX2_30/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3492 OAI22X1_11/a_2_6# INVX2_68/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3493 vdd INVX2_68/Y OAI22X1_11/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3494 gnd INVX2_18/Y OAI22X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3495 OAI22X1_22/a_2_6# INVX2_69/Y OAI22X1_22/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3496 OAI22X1_22/Y OAI22X1_7/D OAI22X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3497 OAI22X1_22/Y INVX2_69/A OAI22X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3498 OAI22X1_22/a_28_54# OAI22X1_7/D OAI22X1_22/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3499 OAI22X1_22/a_9_54# INVX2_18/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3500 OAI22X1_22/a_2_6# INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3501 vdd INVX2_69/Y OAI22X1_22/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3502 DFFNEGX1_7/a_76_6# INVX2_101/Y DFFNEGX1_7/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3503 gnd INVX2_101/Y DFFNEGX1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3504 DFFNEGX1_7/a_66_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3505 INVX2_21/A DFFNEGX1_7/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3506 DFFNEGX1_7/a_23_6# INVX2_101/Y DFFNEGX1_7/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3507 DFFNEGX1_7/a_23_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3508 gnd DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3509 vdd DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3510 DFFNEGX1_7/a_61_74# DFFNEGX1_7/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3511 DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3512 DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3513 vdd INVX2_21/A DFFNEGX1_7/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3514 gnd INVX2_21/A DFFNEGX1_7/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3515 DFFNEGX1_7/a_61_6# DFFNEGX1_7/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3516 DFFNEGX1_7/a_76_84# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3517 INVX2_21/A DFFNEGX1_7/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3518 vdd INVX2_101/Y DFFNEGX1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3519 DFFNEGX1_7/a_31_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3520 DFFNEGX1_7/a_66_6# INVX2_101/Y DFFNEGX1_7/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3521 DFFNEGX1_7/a_17_74# OAI21X1_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3522 DFFNEGX1_7/a_31_74# INVX2_101/Y DFFNEGX1_7/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3523 DFFNEGX1_7/a_17_6# OAI21X1_10/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3524 OAI22X1_8/D NAND2X1_2/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3525 NAND2X1_2/a_9_6# NAND2X1_2/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3526 vdd INVX2_72/Y OAI22X1_8/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3527 OAI22X1_8/D INVX2_72/Y NAND2X1_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3528 INVX2_7/Y INVX2_7/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3529 INVX2_7/Y INVX2_7/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3530 gnd NAND2X1_4/A XNOR2X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3531 NOR2X1_10/A NAND2X1_4/A XNOR2X1_15/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3532 XNOR2X1_15/a_12_41# INVX2_33/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3533 XNOR2X1_15/a_18_54# XNOR2X1_15/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3534 XNOR2X1_15/a_35_6# XNOR2X1_15/a_2_6# NOR2X1_10/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3535 XNOR2X1_15/a_18_6# XNOR2X1_15/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3536 vdd NAND2X1_4/A XNOR2X1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3537 vdd INVX2_33/Y XNOR2X1_15/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3538 NOR2X1_10/A XNOR2X1_15/a_2_6# XNOR2X1_15/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3539 XNOR2X1_15/a_35_54# NAND2X1_4/A NOR2X1_10/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3540 XNOR2X1_15/a_12_41# INVX2_33/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3541 gnd INVX2_33/Y XNOR2X1_15/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3542 gnd INVX2_50/Y XNOR2X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3543 NOR2X1_16/A INVX2_50/Y XNOR2X1_26/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3544 XNOR2X1_26/a_12_41# INVX2_36/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3545 XNOR2X1_26/a_18_54# XNOR2X1_26/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3546 XNOR2X1_26/a_35_6# XNOR2X1_26/a_2_6# NOR2X1_16/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3547 XNOR2X1_26/a_18_6# XNOR2X1_26/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3548 vdd INVX2_50/Y XNOR2X1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3549 vdd INVX2_36/A XNOR2X1_26/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3550 NOR2X1_16/A XNOR2X1_26/a_2_6# XNOR2X1_26/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3551 XNOR2X1_26/a_35_54# INVX2_50/Y NOR2X1_16/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3552 XNOR2X1_26/a_12_41# INVX2_36/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3553 gnd INVX2_36/A XNOR2X1_26/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3554 gnd INVX2_51/Y XNOR2X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3555 NOR2X1_20/B INVX2_51/Y XNOR2X1_37/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3556 XNOR2X1_37/a_12_41# INVX2_28/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3557 XNOR2X1_37/a_18_54# XNOR2X1_37/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3558 XNOR2X1_37/a_35_6# XNOR2X1_37/a_2_6# NOR2X1_20/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3559 XNOR2X1_37/a_18_6# XNOR2X1_37/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3560 vdd INVX2_51/Y XNOR2X1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3561 vdd INVX2_28/A XNOR2X1_37/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3562 NOR2X1_20/B XNOR2X1_37/a_2_6# XNOR2X1_37/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3563 XNOR2X1_37/a_35_54# INVX2_51/Y NOR2X1_20/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3564 XNOR2X1_37/a_12_41# INVX2_28/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3565 gnd INVX2_28/A XNOR2X1_37/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3566 gnd INVX2_57/Y XNOR2X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3567 NOR2X1_27/B INVX2_57/Y XNOR2X1_59/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3568 XNOR2X1_59/a_12_41# INVX2_23/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3569 XNOR2X1_59/a_18_54# XNOR2X1_59/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3570 XNOR2X1_59/a_35_6# XNOR2X1_59/a_2_6# NOR2X1_27/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3571 XNOR2X1_59/a_18_6# XNOR2X1_59/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3572 vdd INVX2_57/Y XNOR2X1_59/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3573 vdd INVX2_23/A XNOR2X1_59/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3574 NOR2X1_27/B XNOR2X1_59/a_2_6# XNOR2X1_59/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3575 XNOR2X1_59/a_35_54# INVX2_57/Y NOR2X1_27/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3576 XNOR2X1_59/a_12_41# INVX2_23/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3577 gnd INVX2_23/A XNOR2X1_59/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3578 gnd INVX2_54/Y XNOR2X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3579 NOR2X1_23/A INVX2_54/Y XNOR2X1_48/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3580 XNOR2X1_48/a_12_41# INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3581 XNOR2X1_48/a_18_54# XNOR2X1_48/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3582 XNOR2X1_48/a_35_6# XNOR2X1_48/a_2_6# NOR2X1_23/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3583 XNOR2X1_48/a_18_6# XNOR2X1_48/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3584 vdd INVX2_54/Y XNOR2X1_48/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3585 vdd INVX2_33/A XNOR2X1_48/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3586 NOR2X1_23/A XNOR2X1_48/a_2_6# XNOR2X1_48/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3587 XNOR2X1_48/a_35_54# INVX2_54/Y NOR2X1_23/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3588 XNOR2X1_48/a_12_41# INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3589 gnd INVX2_33/A XNOR2X1_48/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3590 NOR2X1_5/Y NOR2X1_5/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3591 NOR2X1_5/Y INVX2_1/Y NOR2X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3592 NOR2X1_5/a_9_54# NOR2X1_5/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3593 gnd INVX2_1/Y NOR2X1_5/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3594 gnd INVX2_29/Y OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3595 OAI22X1_12/a_2_6# INVX2_68/Y OAI22X1_12/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3596 OAI22X1_12/Y OAI22X1_9/D OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3597 OAI22X1_12/Y INVX2_68/A OAI22X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3598 OAI22X1_12/a_28_54# OAI22X1_9/D OAI22X1_12/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3599 OAI22X1_12/a_9_54# INVX2_29/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3600 OAI22X1_12/a_2_6# INVX2_68/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3601 vdd INVX2_68/Y OAI22X1_12/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3602 gnd OAI22X1_6/A OAI22X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3603 OAI22X1_23/a_2_6# INVX2_98/Y OAI22X1_23/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3604 OAI22X1_23/Y INVX2_82/Y OAI22X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3605 OAI22X1_23/Y INVX2_57/Y OAI22X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3606 OAI22X1_23/a_28_54# INVX2_82/Y OAI22X1_23/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3607 OAI22X1_23/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3608 OAI22X1_23/a_2_6# INVX2_57/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3609 vdd INVX2_98/Y OAI22X1_23/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3610 DFFNEGX1_8/a_76_6# INVX2_101/Y DFFNEGX1_8/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3611 gnd INVX2_101/Y DFFNEGX1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3612 DFFNEGX1_8/a_66_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3613 NOR2X1_9/B DFFNEGX1_8/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3614 DFFNEGX1_8/a_23_6# INVX2_101/Y DFFNEGX1_8/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3615 DFFNEGX1_8/a_23_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3616 gnd DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3617 vdd DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3618 DFFNEGX1_8/a_61_74# DFFNEGX1_8/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3619 DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3620 DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3621 vdd NOR2X1_9/B DFFNEGX1_8/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3622 gnd NOR2X1_9/B DFFNEGX1_8/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3623 DFFNEGX1_8/a_61_6# DFFNEGX1_8/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3624 DFFNEGX1_8/a_76_84# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3625 NOR2X1_9/B DFFNEGX1_8/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3626 vdd INVX2_101/Y DFFNEGX1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3627 DFFNEGX1_8/a_31_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3628 DFFNEGX1_8/a_66_6# INVX2_101/Y DFFNEGX1_8/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3629 DFFNEGX1_8/a_17_74# OAI21X1_8/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3630 DFFNEGX1_8/a_31_74# INVX2_101/Y DFFNEGX1_8/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3631 DFFNEGX1_8/a_17_6# OAI21X1_8/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3632 OAI22X1_9/D NAND2X1_3/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3633 NAND2X1_3/a_9_6# NAND2X1_3/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3634 vdd INVX2_72/Y OAI22X1_9/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3635 OAI22X1_9/D INVX2_72/Y NAND2X1_3/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3636 INVX2_8/Y INVX2_8/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3637 INVX2_8/Y INVX2_8/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3638 gnd NAND2X1_3/A XNOR2X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3639 NAND3X1_3/B NAND2X1_3/A XNOR2X1_16/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3640 XNOR2X1_16/a_12_41# INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3641 XNOR2X1_16/a_18_54# XNOR2X1_16/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3642 XNOR2X1_16/a_35_6# XNOR2X1_16/a_2_6# NAND3X1_3/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3643 XNOR2X1_16/a_18_6# XNOR2X1_16/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3644 vdd NAND2X1_3/A XNOR2X1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3645 vdd INVX2_32/A XNOR2X1_16/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3646 NAND3X1_3/B XNOR2X1_16/a_2_6# XNOR2X1_16/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3647 XNOR2X1_16/a_35_54# NAND2X1_3/A NAND3X1_3/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3648 XNOR2X1_16/a_12_41# INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3649 gnd INVX2_32/A XNOR2X1_16/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3650 gnd INVX2_50/Y XNOR2X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3651 NOR2X1_20/A INVX2_50/Y XNOR2X1_38/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3652 XNOR2X1_38/a_12_41# INVX2_29/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3653 XNOR2X1_38/a_18_54# XNOR2X1_38/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3654 XNOR2X1_38/a_35_6# XNOR2X1_38/a_2_6# NOR2X1_20/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3655 XNOR2X1_38/a_18_6# XNOR2X1_38/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3656 vdd INVX2_50/Y XNOR2X1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3657 vdd INVX2_29/A XNOR2X1_38/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3658 NOR2X1_20/A XNOR2X1_38/a_2_6# XNOR2X1_38/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3659 XNOR2X1_38/a_35_54# INVX2_50/Y NOR2X1_20/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3660 XNOR2X1_38/a_12_41# INVX2_29/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3661 gnd INVX2_29/A XNOR2X1_38/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3662 gnd INVX2_57/Y XNOR2X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3663 NOR2X1_17/B INVX2_57/Y XNOR2X1_27/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3664 XNOR2X1_27/a_12_41# INVX2_38/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3665 XNOR2X1_27/a_18_54# XNOR2X1_27/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3666 XNOR2X1_27/a_35_6# XNOR2X1_27/a_2_6# NOR2X1_17/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3667 XNOR2X1_27/a_18_6# XNOR2X1_27/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3668 vdd INVX2_57/Y XNOR2X1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3669 vdd INVX2_38/A XNOR2X1_27/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3670 NOR2X1_17/B XNOR2X1_27/a_2_6# XNOR2X1_27/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3671 XNOR2X1_27/a_35_54# INVX2_57/Y NOR2X1_17/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3672 XNOR2X1_27/a_12_41# INVX2_38/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3673 gnd INVX2_38/A XNOR2X1_27/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3674 gnd INVX2_56/Y XNOR2X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3675 NOR2X1_24/B INVX2_56/Y XNOR2X1_49/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3676 XNOR2X1_49/a_12_41# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3677 XNOR2X1_49/a_18_54# XNOR2X1_49/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3678 XNOR2X1_49/a_35_6# XNOR2X1_49/a_2_6# NOR2X1_24/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3679 XNOR2X1_49/a_18_6# XNOR2X1_49/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3680 vdd INVX2_56/Y XNOR2X1_49/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3681 vdd INVX2_31/A XNOR2X1_49/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3682 NOR2X1_24/B XNOR2X1_49/a_2_6# XNOR2X1_49/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3683 XNOR2X1_49/a_35_54# INVX2_56/Y NOR2X1_24/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3684 XNOR2X1_49/a_12_41# INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3685 gnd INVX2_31/A XNOR2X1_49/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3686 NOR2X1_6/Y NOR2X1_6/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3687 NOR2X1_6/Y NOR2X1_6/B NOR2X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3688 NOR2X1_6/a_9_54# NOR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3689 gnd NOR2X1_6/B NOR2X1_6/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3690 gnd INVX2_28/Y OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3691 OAI22X1_13/a_2_6# INVX2_68/Y OAI22X1_13/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3692 OAI22X1_13/Y OAI22X1_8/D OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3693 OAI22X1_13/Y INVX2_68/A OAI22X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3694 OAI22X1_13/a_28_54# OAI22X1_8/D OAI22X1_13/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3695 OAI22X1_13/a_9_54# INVX2_28/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3696 OAI22X1_13/a_2_6# INVX2_68/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3697 vdd INVX2_68/Y OAI22X1_13/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3698 gnd OAI22X1_6/A OAI22X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3699 OAI22X1_24/a_2_6# INVX2_98/Y OAI22X1_24/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3700 OAI22X1_24/Y INVX2_83/Y OAI22X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3701 OAI22X1_24/Y INVX2_56/Y OAI22X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3702 OAI22X1_24/a_28_54# INVX2_83/Y OAI22X1_24/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3703 OAI22X1_24/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3704 OAI22X1_24/a_2_6# INVX2_56/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3705 vdd INVX2_98/Y OAI22X1_24/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3706 DFFNEGX1_9/a_76_6# INVX2_101/Y DFFNEGX1_9/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3707 gnd INVX2_101/Y DFFNEGX1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3708 DFFNEGX1_9/a_66_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3709 INVX2_23/A DFFNEGX1_9/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3710 DFFNEGX1_9/a_23_6# INVX2_101/Y DFFNEGX1_9/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3711 DFFNEGX1_9/a_23_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3712 gnd DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3713 vdd DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3714 DFFNEGX1_9/a_61_74# DFFNEGX1_9/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3715 DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3716 DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3717 vdd INVX2_23/A DFFNEGX1_9/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3718 gnd INVX2_23/A DFFNEGX1_9/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3719 DFFNEGX1_9/a_61_6# DFFNEGX1_9/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3720 DFFNEGX1_9/a_76_84# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3721 INVX2_23/A DFFNEGX1_9/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3722 vdd INVX2_101/Y DFFNEGX1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3723 DFFNEGX1_9/a_31_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3724 DFFNEGX1_9/a_66_6# INVX2_101/Y DFFNEGX1_9/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3725 DFFNEGX1_9/a_17_74# OAI22X1_21/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3726 DFFNEGX1_9/a_31_74# INVX2_101/Y DFFNEGX1_9/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3727 DFFNEGX1_9/a_17_6# OAI22X1_21/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3728 NAND2X1_4/Y NAND2X1_4/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3729 NAND2X1_4/a_9_6# NAND2X1_4/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3730 vdd INVX2_72/Y NAND2X1_4/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3731 NAND2X1_4/Y INVX2_72/Y NAND2X1_4/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3732 INVX2_9/Y INVX2_9/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3733 INVX2_9/Y INVX2_9/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3734 gnd NAND2X1_2/A XNOR2X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3735 NAND3X1_3/A NAND2X1_2/A XNOR2X1_17/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3736 XNOR2X1_17/a_12_41# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3737 XNOR2X1_17/a_18_54# XNOR2X1_17/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3738 XNOR2X1_17/a_35_6# XNOR2X1_17/a_2_6# NAND3X1_3/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3739 XNOR2X1_17/a_18_6# XNOR2X1_17/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3740 vdd NAND2X1_2/A XNOR2X1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3741 vdd INVX2_31/A XNOR2X1_17/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3742 NAND3X1_3/A XNOR2X1_17/a_2_6# XNOR2X1_17/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3743 XNOR2X1_17/a_35_54# NAND2X1_2/A NAND3X1_3/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3744 XNOR2X1_17/a_12_41# INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3745 gnd INVX2_31/A XNOR2X1_17/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3746 gnd INVX2_42/Y XNOR2X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3747 NOR2X1_21/B INVX2_42/Y XNOR2X1_39/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3748 XNOR2X1_39/a_12_41# INVX2_27/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3749 XNOR2X1_39/a_18_54# XNOR2X1_39/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3750 XNOR2X1_39/a_35_6# XNOR2X1_39/a_2_6# NOR2X1_21/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3751 XNOR2X1_39/a_18_6# XNOR2X1_39/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3752 vdd INVX2_42/Y XNOR2X1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3753 vdd INVX2_27/A XNOR2X1_39/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3754 NOR2X1_21/B XNOR2X1_39/a_2_6# XNOR2X1_39/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3755 XNOR2X1_39/a_35_54# INVX2_42/Y NOR2X1_21/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3756 XNOR2X1_39/a_12_41# INVX2_27/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3757 gnd INVX2_27/A XNOR2X1_39/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3758 gnd INVX2_54/Y XNOR2X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3759 NOR2X1_17/A INVX2_54/Y XNOR2X1_28/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3760 XNOR2X1_28/a_12_41# INVX2_35/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3761 XNOR2X1_28/a_18_54# XNOR2X1_28/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3762 XNOR2X1_28/a_35_6# XNOR2X1_28/a_2_6# NOR2X1_17/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3763 XNOR2X1_28/a_18_6# XNOR2X1_28/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3764 vdd INVX2_54/Y XNOR2X1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3765 vdd INVX2_35/A XNOR2X1_28/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3766 NOR2X1_17/A XNOR2X1_28/a_2_6# XNOR2X1_28/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3767 XNOR2X1_28/a_35_54# INVX2_54/Y NOR2X1_17/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3768 XNOR2X1_28/a_12_41# INVX2_35/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3769 gnd INVX2_35/A XNOR2X1_28/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3770 NOR2X1_7/Y NOR2X1_7/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3771 NOR2X1_7/Y NOR2X1_7/B NOR2X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3772 NOR2X1_7/a_9_54# NOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3773 gnd NOR2X1_7/B NOR2X1_7/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3774 gnd INVX2_27/Y OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3775 OAI22X1_14/a_2_6# INVX2_68/Y OAI22X1_14/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3776 OAI22X1_14/Y OAI22X1_7/D OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3777 OAI22X1_14/Y INVX2_68/A OAI22X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3778 OAI22X1_14/a_28_54# OAI22X1_7/D OAI22X1_14/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3779 OAI22X1_14/a_9_54# INVX2_27/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3780 OAI22X1_14/a_2_6# INVX2_68/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3781 vdd INVX2_68/Y OAI22X1_14/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3782 gnd OAI22X1_6/A OAI22X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3783 OAI22X1_25/a_2_6# INVX2_98/Y OAI22X1_25/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3784 OAI22X1_25/Y INVX2_84/Y OAI22X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3785 OAI22X1_25/Y INVX2_55/Y OAI22X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3786 OAI22X1_25/a_28_54# INVX2_84/Y OAI22X1_25/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3787 OAI22X1_25/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3788 OAI22X1_25/a_2_6# INVX2_55/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3789 vdd INVX2_98/Y OAI22X1_25/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3790 OAI21X1_6/B NOR2X1_14/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3791 NAND2X1_5/a_9_6# NOR2X1_14/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3792 vdd NOR2X1_8/B OAI21X1_6/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3793 OAI21X1_6/B NOR2X1_8/B NAND2X1_5/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3794 gnd AOI22X1_3/C XNOR2X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3795 NOR2X1_11/B AOI22X1_3/C XNOR2X1_18/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3796 XNOR2X1_18/a_12_41# INVX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3797 XNOR2X1_18/a_18_54# XNOR2X1_18/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3798 XNOR2X1_18/a_35_6# XNOR2X1_18/a_2_6# NOR2X1_11/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3799 XNOR2X1_18/a_18_6# XNOR2X1_18/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3800 vdd AOI22X1_3/C XNOR2X1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3801 vdd INVX2_23/Y XNOR2X1_18/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3802 NOR2X1_11/B XNOR2X1_18/a_2_6# XNOR2X1_18/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3803 XNOR2X1_18/a_35_54# AOI22X1_3/C NOR2X1_11/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3804 XNOR2X1_18/a_12_41# INVX2_23/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3805 gnd INVX2_23/Y XNOR2X1_18/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3806 gnd INVX2_56/Y XNOR2X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3807 NOR2X1_18/B INVX2_56/Y XNOR2X1_29/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3808 XNOR2X1_29/a_12_41# INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3809 XNOR2X1_29/a_18_54# XNOR2X1_29/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3810 XNOR2X1_29/a_35_6# XNOR2X1_29/a_2_6# NOR2X1_18/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3811 XNOR2X1_29/a_18_6# XNOR2X1_29/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3812 vdd INVX2_56/Y XNOR2X1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3813 vdd INVX2_37/A XNOR2X1_29/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3814 NOR2X1_18/B XNOR2X1_29/a_2_6# XNOR2X1_29/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3815 XNOR2X1_29/a_35_54# INVX2_56/Y NOR2X1_18/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3816 XNOR2X1_29/a_12_41# INVX2_37/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3817 gnd INVX2_37/A XNOR2X1_29/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3818 NOR2X1_8/Y NOR2X1_8/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3819 NOR2X1_8/Y NOR2X1_8/B NOR2X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3820 NOR2X1_8/a_9_54# NOR2X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3821 gnd NOR2X1_8/B NOR2X1_8/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3822 gnd INVX2_33/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3823 OAI22X1_15/a_2_6# INVX2_69/Y OAI22X1_15/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3824 OAI22X1_15/Y NAND2X1_4/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3825 OAI22X1_15/Y INVX2_69/A OAI22X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3826 OAI22X1_15/a_28_54# NAND2X1_4/Y OAI22X1_15/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3827 OAI22X1_15/a_9_54# INVX2_33/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3828 OAI22X1_15/a_2_6# INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3829 vdd INVX2_69/Y OAI22X1_15/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3830 gnd OAI22X1_6/A OAI22X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3831 OAI22X1_26/a_2_6# INVX2_98/Y OAI22X1_26/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3832 OAI22X1_26/Y INVX2_85/Y OAI22X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3833 OAI22X1_26/Y INVX2_54/Y OAI22X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3834 OAI22X1_26/a_28_54# INVX2_85/Y OAI22X1_26/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3835 OAI22X1_26/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3836 OAI22X1_26/a_2_6# INVX2_54/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3837 vdd INVX2_98/Y OAI22X1_26/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3838 OAI21X1_7/C out_valid vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3839 NAND2X1_6/a_9_6# out_valid gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3840 vdd INVX2_65/Y OAI21X1_7/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3841 OAI21X1_7/C INVX2_65/Y NAND2X1_6/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3842 gnd NAND2X1_4/A XNOR2X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3843 NOR2X1_11/A NAND2X1_4/A XNOR2X1_19/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3844 XNOR2X1_19/a_12_41# INVX2_24/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3845 XNOR2X1_19/a_18_54# XNOR2X1_19/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3846 XNOR2X1_19/a_35_6# XNOR2X1_19/a_2_6# NOR2X1_11/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3847 XNOR2X1_19/a_18_6# XNOR2X1_19/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3848 vdd NAND2X1_4/A XNOR2X1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3849 vdd INVX2_24/Y XNOR2X1_19/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3850 NOR2X1_11/A XNOR2X1_19/a_2_6# XNOR2X1_19/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3851 XNOR2X1_19/a_35_54# NAND2X1_4/A NOR2X1_11/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3852 XNOR2X1_19/a_12_41# INVX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3853 gnd INVX2_24/Y XNOR2X1_19/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3854 NOR2X1_9/Y NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3855 NOR2X1_9/Y NOR2X1_9/B NOR2X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3856 NOR2X1_9/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3857 gnd NOR2X1_9/B NOR2X1_9/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3858 gnd INVX2_32/Y OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3859 OAI22X1_16/a_2_6# INVX2_69/Y OAI22X1_16/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3860 OAI22X1_16/Y OAI22X1_9/D OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3861 OAI22X1_16/Y INVX2_69/A OAI22X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3862 OAI22X1_16/a_28_54# OAI22X1_9/D OAI22X1_16/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3863 OAI22X1_16/a_9_54# INVX2_32/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3864 OAI22X1_16/a_2_6# INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3865 vdd INVX2_69/Y OAI22X1_16/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3866 gnd OAI22X1_6/A OAI22X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3867 OAI22X1_27/a_2_6# INVX2_98/Y OAI22X1_27/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3868 OAI22X1_27/Y INVX2_86/Y OAI22X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3869 OAI22X1_27/Y INVX2_52/Y OAI22X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3870 OAI22X1_27/a_28_54# INVX2_86/Y OAI22X1_27/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3871 OAI22X1_27/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3872 OAI22X1_27/a_2_6# INVX2_52/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3873 vdd INVX2_98/Y OAI22X1_27/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3874 NOR2X1_30/Y NOR2X1_30/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3875 NOR2X1_30/Y NOR2X1_30/B NOR2X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3876 NOR2X1_30/a_9_54# NOR2X1_30/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3877 gnd NOR2X1_30/B NOR2X1_30/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3878 OAI21X1_7/B NOR2X1_8/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3879 NAND2X1_7/a_9_6# NOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3880 vdd INVX2_65/A OAI21X1_7/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3881 OAI21X1_7/B INVX2_65/A NAND2X1_7/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3882 gnd INVX2_31/Y OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3883 OAI22X1_17/a_2_6# INVX2_69/Y OAI22X1_17/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3884 OAI22X1_17/Y OAI22X1_8/D OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3885 OAI22X1_17/Y INVX2_69/A OAI22X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3886 OAI22X1_17/a_28_54# OAI22X1_8/D OAI22X1_17/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3887 OAI22X1_17/a_9_54# INVX2_31/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3888 OAI22X1_17/a_2_6# INVX2_69/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3889 vdd INVX2_69/Y OAI22X1_17/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3890 gnd OAI22X1_6/A OAI22X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3891 OAI22X1_28/a_2_6# INVX2_98/Y OAI22X1_28/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3892 OAI22X1_28/Y INVX2_87/Y OAI22X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3893 OAI22X1_28/Y INVX2_51/Y OAI22X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3894 OAI22X1_28/a_28_54# INVX2_87/Y OAI22X1_28/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3895 OAI22X1_28/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3896 OAI22X1_28/a_2_6# INVX2_51/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3897 vdd INVX2_98/Y OAI22X1_28/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3898 NOR2X1_31/Y NOR2X1_31/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3899 NOR2X1_31/Y NOR2X1_31/B NOR2X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3900 NOR2X1_31/a_9_54# NOR2X1_31/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3901 gnd NOR2X1_31/B NOR2X1_31/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3902 NOR2X1_20/Y NOR2X1_20/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3903 NOR2X1_20/Y NOR2X1_20/B NOR2X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3904 NOR2X1_20/a_9_54# NOR2X1_20/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3905 gnd NOR2X1_20/B NOR2X1_20/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3906 NOR2X1_8/A NOR2X1_7/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3907 NAND2X1_8/a_9_6# NOR2X1_7/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3908 vdd NOR2X1_7/A NOR2X1_8/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3909 NOR2X1_8/A NOR2X1_7/A NAND2X1_8/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3910 gnd INVX2_26/Y OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3911 OAI22X1_18/a_2_6# INVX2_71/Y OAI22X1_18/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3912 OAI22X1_18/Y OAI22X1_8/D OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3913 OAI22X1_18/Y INVX2_71/A OAI22X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3914 OAI22X1_18/a_28_54# OAI22X1_8/D OAI22X1_18/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3915 OAI22X1_18/a_9_54# INVX2_26/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3916 OAI22X1_18/a_2_6# INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3917 vdd INVX2_71/Y OAI22X1_18/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3918 gnd OAI22X1_6/A OAI22X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3919 OAI22X1_29/a_2_6# INVX2_98/Y OAI22X1_29/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3920 OAI22X1_29/Y INVX2_88/Y OAI22X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3921 OAI22X1_29/Y INVX2_50/Y OAI22X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3922 OAI22X1_29/a_28_54# INVX2_88/Y OAI22X1_29/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3923 OAI22X1_29/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3924 OAI22X1_29/a_2_6# INVX2_50/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3925 vdd INVX2_98/Y OAI22X1_29/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3926 INVX2_60/A XNOR2X1_82/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M3927 NAND3X1_10/a_9_6# XNOR2X1_82/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M3928 INVX2_60/A NOR2X1_32/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3929 INVX2_60/A NOR2X1_32/Y NAND3X1_10/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M3930 vdd XNOR2X1_81/Y INVX2_60/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3931 NAND3X1_10/a_14_6# XNOR2X1_81/Y NAND3X1_10/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M3932 NOR2X1_10/Y NOR2X1_10/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3933 NOR2X1_10/Y NOR2X1_10/B NOR2X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3934 NOR2X1_10/a_9_54# NOR2X1_10/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3935 gnd NOR2X1_10/B NOR2X1_10/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3936 NOR2X1_21/Y NOR2X1_21/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3937 NOR2X1_21/Y NOR2X1_21/B NOR2X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3938 NOR2X1_21/a_9_54# NOR2X1_21/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3939 gnd NOR2X1_21/B NOR2X1_21/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3940 NOR2X1_32/Y NOR2X1_32/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3941 NOR2X1_32/Y NOR2X1_32/B NOR2X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3942 NOR2X1_32/a_9_54# NOR2X1_32/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3943 gnd NOR2X1_32/B NOR2X1_32/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3944 NAND2X1_9/Y NAND2X1_9/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3945 NAND2X1_9/a_9_6# NAND2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3946 vdd NAND2X1_9/B NAND2X1_9/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3947 NAND2X1_9/Y NAND2X1_9/B NAND2X1_9/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3948 gnd INVX2_25/Y OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3949 OAI22X1_19/a_2_6# INVX2_71/Y OAI22X1_19/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3950 OAI22X1_19/Y OAI22X1_9/D OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3951 OAI22X1_19/Y INVX2_71/A OAI22X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3952 OAI22X1_19/a_28_54# OAI22X1_9/D OAI22X1_19/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3953 OAI22X1_19/a_9_54# INVX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3954 OAI22X1_19/a_2_6# INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3955 vdd INVX2_71/Y OAI22X1_19/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3956 INVX2_48/A XNOR2X1_86/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M3957 NAND3X1_11/a_9_6# XNOR2X1_86/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M3958 INVX2_48/A NOR2X1_33/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3959 INVX2_48/A NOR2X1_33/Y NAND3X1_11/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M3960 vdd XNOR2X1_85/Y INVX2_48/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3961 NAND3X1_11/a_14_6# XNOR2X1_85/Y NAND3X1_11/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M3962 NOR2X1_11/Y NOR2X1_11/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3963 NOR2X1_11/Y NOR2X1_11/B NOR2X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3964 NOR2X1_11/a_9_54# NOR2X1_11/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3965 gnd NOR2X1_11/B NOR2X1_11/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3966 NOR2X1_33/Y NOR2X1_33/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3967 NOR2X1_33/Y NOR2X1_33/B NOR2X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3968 NOR2X1_33/a_9_54# NOR2X1_33/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3969 gnd NOR2X1_33/B NOR2X1_33/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3970 NOR2X1_22/Y NOR2X1_22/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3971 NOR2X1_22/Y NOR2X1_22/B NOR2X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3972 NOR2X1_22/a_9_54# NOR2X1_22/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3973 gnd NOR2X1_22/B NOR2X1_22/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3974 INVX2_90/Y in_ans0[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3975 INVX2_90/Y in_ans0[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3976 gnd OAI21X1_20/A OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3977 vdd AOI22X1_8/Y XOR2X1_4/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3978 XOR2X1_4/A AOI22X1_8/Y OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3979 XOR2X1_4/A OAI21X1_20/B OAI21X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3980 OAI21X1_20/a_9_54# OAI21X1_20/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3981 OAI21X1_20/a_2_6# OAI21X1_20/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3982 INVX2_70/A NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3983 INVX2_70/A OR2X1_0/B NOR2X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3984 NOR2X1_12/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3985 gnd OR2X1_0/B INVX2_70/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3986 INVX2_43/A XNOR2X1_90/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M3987 NAND3X1_12/a_9_6# XNOR2X1_90/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M3988 INVX2_43/A NOR2X1_34/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3989 INVX2_43/A NOR2X1_34/Y NAND3X1_12/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M3990 vdd XNOR2X1_89/Y INVX2_43/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3991 NAND3X1_12/a_14_6# XNOR2X1_89/Y NAND3X1_12/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M3992 NOR2X1_34/Y NOR2X1_34/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3993 NOR2X1_34/Y NOR2X1_34/B NOR2X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3994 NOR2X1_34/a_9_54# NOR2X1_34/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3995 gnd NOR2X1_34/B NOR2X1_34/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3996 NOR2X1_23/Y NOR2X1_23/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M3997 NOR2X1_23/Y NOR2X1_23/B NOR2X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M3998 NOR2X1_23/a_9_54# NOR2X1_23/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3999 gnd NOR2X1_23/B NOR2X1_23/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4000 DFFSR_0/a_23_27# DFFSR_0/a_47_71# DFFSR_0/a_2_6# vdd pfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M4001 DFFSR_0/a_2_6# DFFSR_0/R vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M4002 DFFSR_0/a_47_71# BUFX2_0/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M4003 DFFSR_0/a_47_71# BUFX2_0/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M4004 DFFSR_0/a_113_6# DFFSR_7/S DFFSR_0/a_146_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=40p ps=24u
M4005 DFFSR_0/a_10_61# DFFSR_0/a_23_27# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M4006 DFFSR_0/a_113_6# DFFSR_0/a_47_4# DFFSR_0/a_105_6# vdd pfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M4007 vdd DFFSR_0/a_122_6# DFFSR_1/D vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M4008 vdd DFFSR_7/S DFFSR_0/a_113_6# vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M4009 DFFSR_0/a_26_6# DFFSR_0/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=40p pd=24u as=80p ps=28u
M4010 DFFSR_0/a_23_27# DFFSR_0/a_47_4# DFFSR_0/a_2_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M4011 DFFSR_0/a_57_6# DFFSR_0/a_47_4# DFFSR_0/a_23_27# vdd pfet w=10 l=2
+  ad=55p pd=26u as=29.999998p ps=16u
M4012 gnd DFFSR_0/a_10_61# DFFSR_0/a_10_6# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=40p ps=24u
M4013 DFFSR_0/a_105_6# DFFSR_0/a_47_4# DFFSR_0/a_10_61# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M4014 vdd DFFSR_7/S DFFSR_0/a_10_61# vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M4015 gnd DFFSR_0/D DFFSR_0/a_57_6# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M4016 DFFSR_0/a_122_6# DFFSR_0/a_105_6# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M4017 DFFSR_0/a_10_61# DFFSR_7/S DFFSR_0/a_26_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=40p ps=24u
M4018 gnd DFFSR_0/a_47_71# DFFSR_0/a_47_4# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M4019 vdd DFFSR_0/R DFFSR_0/a_122_6# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M4020 DFFSR_0/a_130_6# DFFSR_0/a_105_6# DFFSR_0/a_122_6# Gnd nfet w=20 l=2
+  ad=40p pd=24u as=0.12n ps=52u
M4021 DFFSR_0/a_10_6# DFFSR_0/R DFFSR_0/a_2_6# Gnd nfet w=20 l=2
+  ad=40p pd=24u as=0.12n ps=52u
M4022 vdd DFFSR_0/a_47_71# DFFSR_0/a_47_4# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M4023 DFFSR_0/a_57_6# DFFSR_0/a_47_71# DFFSR_0/a_23_27# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=29.999998p ps=16u
M4024 vdd DFFSR_0/D DFFSR_0/a_57_6# vdd pfet w=20 l=2
+  ad=100p pd=50u as=55p ps=26u
M4025 vdd DFFSR_0/a_10_61# DFFSR_0/a_2_6# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M4026 DFFSR_0/a_105_6# DFFSR_0/a_47_71# DFFSR_0/a_10_61# vdd pfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M4027 DFFSR_0/a_146_6# DFFSR_0/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=40p pd=24u as=80p ps=28u
M4028 gnd DFFSR_0/a_122_6# DFFSR_1/D Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M4029 DFFSR_0/a_113_6# DFFSR_0/a_122_6# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M4030 DFFSR_0/a_113_6# DFFSR_0/a_47_71# DFFSR_0/a_105_6# Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M4031 gnd DFFSR_0/R DFFSR_0/a_130_6# Gnd nfet w=20 l=2
+  ad=80p pd=28u as=40p ps=24u
M4032 INVX2_80/Y in_ans3[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4033 INVX2_80/Y in_ans3[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4034 INVX2_91/Y in_ans0[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4035 INVX2_91/Y in_ans0[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4036 gnd in_loadtest OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4037 vdd OAI21X1_21/C OAI21X1_21/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4038 OAI21X1_21/Y OAI21X1_21/C OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4039 OAI21X1_21/Y INVX2_63/Y OAI21X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4040 OAI21X1_21/a_9_54# in_loadtest vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4041 OAI21X1_21/a_2_6# INVX2_63/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4042 gnd NOR2X1_6/A OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4043 vdd NAND3X1_2/Y OAI21X1_10/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4044 OAI21X1_10/Y NAND3X1_2/Y OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4045 OAI21X1_10/Y NOR2X1_7/B OAI21X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4046 OAI21X1_10/a_9_54# NOR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4047 OAI21X1_10/a_2_6# NOR2X1_7/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4048 NOR2X1_35/Y INVX2_62/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4049 NOR2X1_35/Y out_state[1] NOR2X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4050 NOR2X1_35/a_9_54# INVX2_62/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4051 gnd out_state[1] NOR2X1_35/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4052 NOR2X1_13/Y INVX2_99/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4053 NOR2X1_13/Y OR2X1_0/B NOR2X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4054 NOR2X1_13/a_9_54# INVX2_99/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4055 gnd OR2X1_0/B NOR2X1_13/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4056 NOR2X1_24/Y NOR2X1_24/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4057 NOR2X1_24/Y NOR2X1_24/B NOR2X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4058 NOR2X1_24/a_9_54# NOR2X1_24/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4059 gnd NOR2X1_24/B NOR2X1_24/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4060 DFFSR_1/a_23_27# DFFSR_1/a_47_71# DFFSR_1/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4061 DFFSR_1/a_2_6# DFFSR_1/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4062 DFFSR_1/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4063 DFFSR_1/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4064 DFFSR_1/a_113_6# DFFSR_7/S DFFSR_1/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4065 DFFSR_1/a_10_61# DFFSR_1/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4066 DFFSR_1/a_113_6# DFFSR_1/a_47_4# DFFSR_1/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4067 vdd DFFSR_1/a_122_6# DFFSR_2/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4068 vdd DFFSR_7/S DFFSR_1/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4069 DFFSR_1/a_26_6# DFFSR_1/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4070 DFFSR_1/a_23_27# DFFSR_1/a_47_4# DFFSR_1/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4071 DFFSR_1/a_57_6# DFFSR_1/a_47_4# DFFSR_1/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4072 gnd DFFSR_1/a_10_61# DFFSR_1/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4073 DFFSR_1/a_105_6# DFFSR_1/a_47_4# DFFSR_1/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4074 vdd DFFSR_7/S DFFSR_1/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4075 gnd DFFSR_1/D DFFSR_1/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4076 DFFSR_1/a_122_6# DFFSR_1/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4077 DFFSR_1/a_10_61# DFFSR_7/S DFFSR_1/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4078 gnd DFFSR_1/a_47_71# DFFSR_1/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4079 vdd DFFSR_1/R DFFSR_1/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4080 DFFSR_1/a_130_6# DFFSR_1/a_105_6# DFFSR_1/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4081 DFFSR_1/a_10_6# DFFSR_1/R DFFSR_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4082 vdd DFFSR_1/a_47_71# DFFSR_1/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4083 DFFSR_1/a_57_6# DFFSR_1/a_47_71# DFFSR_1/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4084 vdd DFFSR_1/D DFFSR_1/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4085 vdd DFFSR_1/a_10_61# DFFSR_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4086 DFFSR_1/a_105_6# DFFSR_1/a_47_71# DFFSR_1/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4087 DFFSR_1/a_146_6# DFFSR_1/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4088 gnd DFFSR_1/a_122_6# DFFSR_2/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4089 DFFSR_1/a_113_6# DFFSR_1/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4090 DFFSR_1/a_113_6# DFFSR_1/a_47_71# DFFSR_1/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4091 gnd DFFSR_1/R DFFSR_1/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4092 INVX2_70/Y INVX2_70/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4093 INVX2_70/Y INVX2_70/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4094 INVX2_92/Y in_ans0[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4095 INVX2_92/Y in_ans0[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4096 INVX2_81/Y in_ans3[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4097 INVX2_81/Y in_ans3[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4098 gnd AOI21X1_2/Y OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4099 vdd OAI21X1_12/Y INVX2_73/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4100 INVX2_73/A OAI21X1_12/Y OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4101 INVX2_73/A INVX2_65/A OAI21X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4102 OAI21X1_11/a_9_54# AOI21X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4103 OAI21X1_11/a_2_6# INVX2_65/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4104 gnd out_state[1] OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4105 vdd INVX2_62/Y AND2X2_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4106 AND2X2_4/B INVX2_62/Y OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4107 AND2X2_4/B INVX2_95/Y OAI21X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4108 OAI21X1_22/a_9_54# out_state[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4109 OAI21X1_22/a_2_6# INVX2_95/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4110 NOR2X1_36/Y INVX2_63/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4111 NOR2X1_36/Y INVX2_62/Y NOR2X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4112 NOR2X1_36/a_9_54# INVX2_63/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4113 gnd INVX2_62/Y NOR2X1_36/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4114 NOR2X1_14/Y NOR2X1_7/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4115 NOR2X1_14/Y INVX2_21/A NOR2X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4116 NOR2X1_14/a_9_54# NOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4117 gnd INVX2_21/A NOR2X1_14/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4118 NOR2X1_25/Y NOR2X1_25/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4119 NOR2X1_25/Y NOR2X1_25/B NOR2X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4120 NOR2X1_25/a_9_54# NOR2X1_25/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4121 gnd NOR2X1_25/B NOR2X1_25/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4122 gnd INVX2_7/A MUX2X1_10/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4123 MUX2X1_10/a_17_50# INVX2_7/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4124 INVX2_9/A MUX2X1_9/S MUX2X1_10/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4125 MUX2X1_10/a_30_54# MUX2X1_10/a_2_10# INVX2_9/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4126 MUX2X1_10/a_17_10# INVX2_7/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4127 vdd MUX2X1_9/S MUX2X1_10/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4128 MUX2X1_10/a_30_10# MUX2X1_9/S INVX2_9/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4129 gnd MUX2X1_9/S MUX2X1_10/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4130 vdd INVX2_7/A MUX2X1_10/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4131 INVX2_9/A MUX2X1_10/a_2_10# MUX2X1_10/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4132 DFFSR_2/a_23_27# DFFSR_2/a_47_71# DFFSR_2/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4133 DFFSR_2/a_2_6# DFFSR_2/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4134 DFFSR_2/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4135 DFFSR_2/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4136 DFFSR_2/a_113_6# DFFSR_7/S DFFSR_2/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4137 DFFSR_2/a_10_61# DFFSR_2/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4138 DFFSR_2/a_113_6# DFFSR_2/a_47_4# DFFSR_2/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4139 vdd DFFSR_2/a_122_6# DFFSR_3/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4140 vdd DFFSR_7/S DFFSR_2/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4141 DFFSR_2/a_26_6# DFFSR_2/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4142 DFFSR_2/a_23_27# DFFSR_2/a_47_4# DFFSR_2/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4143 DFFSR_2/a_57_6# DFFSR_2/a_47_4# DFFSR_2/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4144 gnd DFFSR_2/a_10_61# DFFSR_2/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4145 DFFSR_2/a_105_6# DFFSR_2/a_47_4# DFFSR_2/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4146 vdd DFFSR_7/S DFFSR_2/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4147 gnd DFFSR_2/D DFFSR_2/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4148 DFFSR_2/a_122_6# DFFSR_2/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4149 DFFSR_2/a_10_61# DFFSR_7/S DFFSR_2/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4150 gnd DFFSR_2/a_47_71# DFFSR_2/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4151 vdd DFFSR_2/R DFFSR_2/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4152 DFFSR_2/a_130_6# DFFSR_2/a_105_6# DFFSR_2/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4153 DFFSR_2/a_10_6# DFFSR_2/R DFFSR_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4154 vdd DFFSR_2/a_47_71# DFFSR_2/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4155 DFFSR_2/a_57_6# DFFSR_2/a_47_71# DFFSR_2/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4156 vdd DFFSR_2/D DFFSR_2/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4157 vdd DFFSR_2/a_10_61# DFFSR_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4158 DFFSR_2/a_105_6# DFFSR_2/a_47_71# DFFSR_2/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4159 DFFSR_2/a_146_6# DFFSR_2/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4160 gnd DFFSR_2/a_122_6# DFFSR_3/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4161 DFFSR_2/a_113_6# DFFSR_2/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4162 DFFSR_2/a_113_6# DFFSR_2/a_47_71# DFFSR_2/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4163 gnd DFFSR_2/R DFFSR_2/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4164 INVX2_71/Y INVX2_71/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4165 INVX2_71/Y INVX2_71/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4166 INVX2_82/Y in_ans2[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4167 INVX2_82/Y in_ans2[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4168 INVX2_93/Y in_ans0[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4169 INVX2_93/Y in_ans0[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4170 INVX2_60/Y INVX2_60/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4171 INVX2_60/Y INVX2_60/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4172 gnd OR2X1_0/B OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4173 vdd INVX2_72/Y OAI21X1_12/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4174 OAI21X1_12/Y INVX2_72/Y OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4175 OAI21X1_12/Y OR2X1_0/A OAI21X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4176 OAI21X1_12/a_9_54# OR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4177 OAI21X1_12/a_2_6# OR2X1_0/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4178 NOR2X1_37/Y in_restart gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4179 NOR2X1_37/Y NOR2X1_37/B NOR2X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4180 NOR2X1_37/a_9_54# in_restart vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4181 gnd NOR2X1_37/B NOR2X1_37/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4182 NOR2X1_15/Y NOR2X1_15/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4183 NOR2X1_15/Y NOR2X1_15/B NOR2X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4184 NOR2X1_15/a_9_54# NOR2X1_15/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4185 gnd NOR2X1_15/B NOR2X1_15/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4186 NOR2X1_26/Y NOR2X1_26/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4187 NOR2X1_26/Y NOR2X1_26/B NOR2X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4188 NOR2X1_26/a_9_54# NOR2X1_26/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4189 gnd NOR2X1_26/B NOR2X1_26/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4190 gnd DFFSR_3/D MUX2X1_11/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4191 MUX2X1_11/a_17_50# DFFSR_3/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4192 INVX2_10/A MUX2X1_9/S MUX2X1_11/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4193 MUX2X1_11/a_30_54# MUX2X1_11/a_2_10# INVX2_10/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4194 MUX2X1_11/a_17_10# DFFSR_3/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4195 vdd MUX2X1_9/S MUX2X1_11/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4196 MUX2X1_11/a_30_10# MUX2X1_9/S INVX2_10/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4197 gnd MUX2X1_9/S MUX2X1_11/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4198 vdd DFFSR_3/D MUX2X1_11/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4199 INVX2_10/A MUX2X1_11/a_2_10# MUX2X1_11/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4200 DFFSR_3/a_23_27# DFFSR_3/a_47_71# DFFSR_3/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4201 DFFSR_3/a_2_6# DFFSR_3/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4202 DFFSR_3/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4203 DFFSR_3/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4204 DFFSR_3/a_113_6# DFFSR_7/S DFFSR_3/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4205 DFFSR_3/a_10_61# DFFSR_3/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4206 DFFSR_3/a_113_6# DFFSR_3/a_47_4# DFFSR_3/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4207 vdd DFFSR_3/a_122_6# DFFSR_4/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4208 vdd DFFSR_7/S DFFSR_3/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4209 DFFSR_3/a_26_6# DFFSR_3/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4210 DFFSR_3/a_23_27# DFFSR_3/a_47_4# DFFSR_3/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4211 DFFSR_3/a_57_6# DFFSR_3/a_47_4# DFFSR_3/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4212 gnd DFFSR_3/a_10_61# DFFSR_3/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4213 DFFSR_3/a_105_6# DFFSR_3/a_47_4# DFFSR_3/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4214 vdd DFFSR_7/S DFFSR_3/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4215 gnd DFFSR_3/D DFFSR_3/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4216 DFFSR_3/a_122_6# DFFSR_3/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4217 DFFSR_3/a_10_61# DFFSR_7/S DFFSR_3/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4218 gnd DFFSR_3/a_47_71# DFFSR_3/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4219 vdd DFFSR_3/R DFFSR_3/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4220 DFFSR_3/a_130_6# DFFSR_3/a_105_6# DFFSR_3/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4221 DFFSR_3/a_10_6# DFFSR_3/R DFFSR_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4222 vdd DFFSR_3/a_47_71# DFFSR_3/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4223 DFFSR_3/a_57_6# DFFSR_3/a_47_71# DFFSR_3/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4224 vdd DFFSR_3/D DFFSR_3/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4225 vdd DFFSR_3/a_10_61# DFFSR_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4226 DFFSR_3/a_105_6# DFFSR_3/a_47_71# DFFSR_3/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4227 DFFSR_3/a_146_6# DFFSR_3/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4228 gnd DFFSR_3/a_122_6# DFFSR_4/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4229 DFFSR_3/a_113_6# DFFSR_3/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4230 DFFSR_3/a_113_6# DFFSR_3/a_47_71# DFFSR_3/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4231 gnd DFFSR_3/R DFFSR_3/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4232 INVX2_94/Y in_restart gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4233 INVX2_94/Y in_restart vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4234 INVX2_72/Y NOR2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4235 INVX2_72/Y NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4236 INVX2_50/Y INVX2_50/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4237 INVX2_50/Y INVX2_50/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4238 out_Anum[2] INVX2_61/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4239 out_Anum[2] INVX2_61/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4240 INVX2_83/Y in_ans2[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4241 INVX2_83/Y in_ans2[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4242 gnd AOI21X1_1/Y OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4243 vdd DFFSR_7/S INVX2_65/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4244 INVX2_65/A DFFSR_7/S OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4245 INVX2_65/A NOR2X1_9/A OAI21X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4246 OAI21X1_13/a_9_54# AOI21X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4247 OAI21X1_13/a_2_6# NOR2X1_9/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4248 gnd NOR2X1_0/B XNOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4249 XNOR2X1_0/Y NOR2X1_0/B XNOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4250 XNOR2X1_0/a_12_41# NOR2X1_0/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4251 XNOR2X1_0/a_18_54# XNOR2X1_0/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4252 XNOR2X1_0/a_35_6# XNOR2X1_0/a_2_6# XNOR2X1_0/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4253 XNOR2X1_0/a_18_6# XNOR2X1_0/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4254 vdd NOR2X1_0/B XNOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4255 vdd NOR2X1_0/A XNOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4256 XNOR2X1_0/Y XNOR2X1_0/a_2_6# XNOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4257 XNOR2X1_0/a_35_54# NOR2X1_0/B XNOR2X1_0/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4258 XNOR2X1_0/a_12_41# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4259 gnd NOR2X1_0/A XNOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4260 INVX4_0/A in_clkb vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M4261 INVX4_0/A in_clkb gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M4262 AND2X2_0/a_2_6# DFFSR_7/S vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M4263 AND2X2_0/a_9_6# DFFSR_7/S AND2X2_0/a_2_6# Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M4264 AND2X2_0/Y AND2X2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M4265 AND2X2_0/Y AND2X2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.108n ps=46u
M4266 vdd INVX2_98/Y AND2X2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0.108n pd=46u as=59.999996p ps=26u
M4267 gnd INVX2_98/Y AND2X2_0/a_9_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=29.999998p ps=23u
M4268 NOR2X1_16/Y NOR2X1_16/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4269 NOR2X1_16/Y NOR2X1_16/B NOR2X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4270 NOR2X1_16/a_9_54# NOR2X1_16/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4271 gnd NOR2X1_16/B NOR2X1_16/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4272 NOR2X1_27/Y NOR2X1_27/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4273 NOR2X1_27/Y NOR2X1_27/B NOR2X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4274 NOR2X1_27/a_9_54# NOR2X1_27/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4275 gnd NOR2X1_27/B NOR2X1_27/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4276 gnd XNOR2X1_3/Y MUX2X1_12/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4277 MUX2X1_12/a_17_50# INVX2_8/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4278 OAI21X1_0/C OAI21X1_1/Y MUX2X1_12/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4279 MUX2X1_12/a_30_54# MUX2X1_12/a_2_10# OAI21X1_0/C vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4280 MUX2X1_12/a_17_10# INVX2_8/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4281 vdd OAI21X1_1/Y MUX2X1_12/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4282 MUX2X1_12/a_30_10# OAI21X1_1/Y OAI21X1_0/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4283 gnd OAI21X1_1/Y MUX2X1_12/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4284 vdd XNOR2X1_3/Y MUX2X1_12/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4285 OAI21X1_0/C MUX2X1_12/a_2_10# MUX2X1_12/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4286 DFFSR_4/a_23_27# DFFSR_4/a_47_71# DFFSR_4/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4287 DFFSR_4/a_2_6# DFFSR_4/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4288 DFFSR_4/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4289 DFFSR_4/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4290 DFFSR_4/a_113_6# DFFSR_7/S DFFSR_4/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4291 DFFSR_4/a_10_61# DFFSR_4/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4292 DFFSR_4/a_113_6# DFFSR_4/a_47_4# DFFSR_4/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4293 vdd DFFSR_4/a_122_6# DFFSR_5/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4294 vdd DFFSR_7/S DFFSR_4/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4295 DFFSR_4/a_26_6# DFFSR_4/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4296 DFFSR_4/a_23_27# DFFSR_4/a_47_4# DFFSR_4/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4297 DFFSR_4/a_57_6# DFFSR_4/a_47_4# DFFSR_4/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4298 gnd DFFSR_4/a_10_61# DFFSR_4/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4299 DFFSR_4/a_105_6# DFFSR_4/a_47_4# DFFSR_4/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4300 vdd DFFSR_7/S DFFSR_4/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4301 gnd DFFSR_4/D DFFSR_4/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4302 DFFSR_4/a_122_6# DFFSR_4/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4303 DFFSR_4/a_10_61# DFFSR_7/S DFFSR_4/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4304 gnd DFFSR_4/a_47_71# DFFSR_4/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4305 vdd DFFSR_4/R DFFSR_4/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4306 DFFSR_4/a_130_6# DFFSR_4/a_105_6# DFFSR_4/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4307 DFFSR_4/a_10_6# DFFSR_4/R DFFSR_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4308 vdd DFFSR_4/a_47_71# DFFSR_4/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4309 DFFSR_4/a_57_6# DFFSR_4/a_47_71# DFFSR_4/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4310 vdd DFFSR_4/D DFFSR_4/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4311 vdd DFFSR_4/a_10_61# DFFSR_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4312 DFFSR_4/a_105_6# DFFSR_4/a_47_71# DFFSR_4/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4313 DFFSR_4/a_146_6# DFFSR_4/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4314 gnd DFFSR_4/a_122_6# DFFSR_5/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4315 DFFSR_4/a_113_6# DFFSR_4/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4316 DFFSR_4/a_113_6# DFFSR_4/a_47_71# DFFSR_4/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4317 gnd DFFSR_4/R DFFSR_4/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4318 INVX2_62/Y out_state[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4319 INVX2_62/Y out_state[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4320 INVX2_73/Y INVX2_73/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4321 INVX2_73/Y INVX2_73/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4322 INVX2_51/Y INVX2_51/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4323 INVX2_51/Y INVX2_51/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4324 INVX2_40/Y INVX2_40/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4325 INVX2_40/Y INVX2_40/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4326 INVX2_95/Y in_loadtest gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4327 INVX2_95/Y in_loadtest vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4328 INVX2_84/Y in_ans2[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4329 INVX2_84/Y in_ans2[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4330 gnd OAI21X1_14/A OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4331 vdd AND2X2_2/Y INVX2_34/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4332 INVX2_34/A AND2X2_2/Y OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4333 INVX2_34/A NAND2X1_9/Y OAI21X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4334 OAI21X1_14/a_9_54# OAI21X1_14/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4335 OAI21X1_14/a_2_6# NAND2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4336 gnd INVX2_11/Y XNOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4337 XNOR2X1_1/Y INVX2_11/Y XNOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4338 XNOR2X1_1/a_12_41# NOR2X1_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4339 XNOR2X1_1/a_18_54# XNOR2X1_1/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4340 XNOR2X1_1/a_35_6# XNOR2X1_1/a_2_6# XNOR2X1_1/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4341 XNOR2X1_1/a_18_6# XNOR2X1_1/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4342 vdd INVX2_11/Y XNOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4343 vdd NOR2X1_0/Y XNOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4344 XNOR2X1_1/Y XNOR2X1_1/a_2_6# XNOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4345 XNOR2X1_1/a_35_54# INVX2_11/Y XNOR2X1_1/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4346 XNOR2X1_1/a_12_41# NOR2X1_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4347 gnd NOR2X1_0/Y XNOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4348 AND2X2_1/a_2_6# NOR2X1_9/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4349 AND2X2_1/a_9_6# NOR2X1_9/B AND2X2_1/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M4350 OR2X1_0/A AND2X2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4351 OR2X1_0/A AND2X2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4352 vdd NOR2X1_8/A AND2X2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4353 gnd NOR2X1_8/A AND2X2_1/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4354 NOR2X1_28/Y NOR2X1_28/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4355 NOR2X1_28/Y NOR2X1_28/B NOR2X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4356 NOR2X1_28/a_9_54# NOR2X1_28/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4357 gnd NOR2X1_28/B NOR2X1_28/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4358 NOR2X1_17/Y NOR2X1_17/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4359 NOR2X1_17/Y NOR2X1_17/B NOR2X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4360 NOR2X1_17/a_9_54# NOR2X1_17/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4361 gnd NOR2X1_17/B NOR2X1_17/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4362 gnd XNOR2X1_2/Y MUX2X1_13/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4363 MUX2X1_13/a_17_50# INVX2_9/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4364 INVX2_11/A OAI21X1_1/Y MUX2X1_13/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4365 MUX2X1_13/a_30_54# MUX2X1_13/a_2_10# INVX2_11/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4366 MUX2X1_13/a_17_10# INVX2_9/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4367 vdd OAI21X1_1/Y MUX2X1_13/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4368 MUX2X1_13/a_30_10# OAI21X1_1/Y INVX2_11/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4369 gnd OAI21X1_1/Y MUX2X1_13/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4370 vdd XNOR2X1_2/Y MUX2X1_13/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4371 INVX2_11/A MUX2X1_13/a_2_10# MUX2X1_13/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4372 DFFSR_5/a_23_27# DFFSR_5/a_47_71# DFFSR_5/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4373 DFFSR_5/a_2_6# DFFSR_5/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4374 DFFSR_5/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4375 DFFSR_5/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4376 DFFSR_5/a_113_6# DFFSR_7/S DFFSR_5/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4377 DFFSR_5/a_10_61# DFFSR_5/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4378 DFFSR_5/a_113_6# DFFSR_5/a_47_4# DFFSR_5/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4379 vdd DFFSR_5/a_122_6# INVX2_0/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4380 vdd DFFSR_7/S DFFSR_5/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4381 DFFSR_5/a_26_6# DFFSR_5/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4382 DFFSR_5/a_23_27# DFFSR_5/a_47_4# DFFSR_5/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4383 DFFSR_5/a_57_6# DFFSR_5/a_47_4# DFFSR_5/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4384 gnd DFFSR_5/a_10_61# DFFSR_5/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4385 DFFSR_5/a_105_6# DFFSR_5/a_47_4# DFFSR_5/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4386 vdd DFFSR_7/S DFFSR_5/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4387 gnd DFFSR_5/D DFFSR_5/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4388 DFFSR_5/a_122_6# DFFSR_5/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4389 DFFSR_5/a_10_61# DFFSR_7/S DFFSR_5/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4390 gnd DFFSR_5/a_47_71# DFFSR_5/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4391 vdd DFFSR_5/R DFFSR_5/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4392 DFFSR_5/a_130_6# DFFSR_5/a_105_6# DFFSR_5/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4393 DFFSR_5/a_10_6# DFFSR_5/R DFFSR_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4394 vdd DFFSR_5/a_47_71# DFFSR_5/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4395 DFFSR_5/a_57_6# DFFSR_5/a_47_71# DFFSR_5/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4396 vdd DFFSR_5/D DFFSR_5/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4397 vdd DFFSR_5/a_10_61# DFFSR_5/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4398 DFFSR_5/a_105_6# DFFSR_5/a_47_71# DFFSR_5/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4399 DFFSR_5/a_146_6# DFFSR_5/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4400 gnd DFFSR_5/a_122_6# INVX2_0/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4401 DFFSR_5/a_113_6# DFFSR_5/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4402 DFFSR_5/a_113_6# DFFSR_5/a_47_71# DFFSR_5/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4403 gnd DFFSR_5/R DFFSR_5/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4404 INVX2_63/Y out_state[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4405 INVX2_63/Y out_state[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4406 BUFX2_1/A in_clka gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4407 BUFX2_1/A in_clka vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4408 INVX2_74/Y INVX2_74/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4409 INVX2_74/Y INVX2_74/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4410 INVX2_30/Y INVX2_30/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4411 INVX2_30/Y INVX2_30/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4412 INVX2_85/Y in_ans2[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4413 INVX2_85/Y in_ans2[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4414 INVX2_52/Y INVX2_52/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4415 INVX2_52/Y INVX2_52/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4416 INVX2_41/Y INVX2_41/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4417 INVX2_41/Y INVX2_41/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4418 gnd NOR2X1_7/A OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4419 vdd AND2X2_3/B AOI21X1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4420 AOI21X1_2/B AND2X2_3/B OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4421 AOI21X1_2/B AND2X2_2/B OAI21X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4422 OAI21X1_15/a_9_54# NOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4423 OAI21X1_15/a_2_6# AND2X2_2/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4424 gnd NOR2X1_1/B XNOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4425 XNOR2X1_2/Y NOR2X1_1/B XNOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4426 XNOR2X1_2/a_12_41# INVX2_9/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4427 XNOR2X1_2/a_18_54# XNOR2X1_2/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4428 XNOR2X1_2/a_35_6# XNOR2X1_2/a_2_6# XNOR2X1_2/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4429 XNOR2X1_2/a_18_6# XNOR2X1_2/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4430 vdd NOR2X1_1/B XNOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4431 vdd INVX2_9/Y XNOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4432 XNOR2X1_2/Y XNOR2X1_2/a_2_6# XNOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4433 XNOR2X1_2/a_35_54# NOR2X1_1/B XNOR2X1_2/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4434 XNOR2X1_2/a_12_41# INVX2_9/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4435 gnd INVX2_9/Y XNOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4436 AND2X2_2/a_2_6# AND2X2_3/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4437 AND2X2_2/a_9_6# AND2X2_3/B AND2X2_2/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M4438 AND2X2_2/Y AND2X2_2/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4439 AND2X2_2/Y AND2X2_2/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4440 vdd AND2X2_2/B AND2X2_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4441 gnd AND2X2_2/B AND2X2_2/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4442 NOR2X1_29/Y NOR2X1_29/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4443 NOR2X1_29/Y NOR2X1_29/B NOR2X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4444 NOR2X1_29/a_9_54# NOR2X1_29/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4445 gnd NOR2X1_29/B NOR2X1_29/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4446 NOR2X1_18/Y NOR2X1_18/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4447 NOR2X1_18/Y NOR2X1_18/B NOR2X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4448 NOR2X1_18/a_9_54# NOR2X1_18/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4449 gnd NOR2X1_18/B NOR2X1_18/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4450 gnd INVX2_10/A MUX2X1_14/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4451 MUX2X1_14/a_17_50# NOR2X1_1/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4452 INVX2_12/A OAI21X1_1/Y MUX2X1_14/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4453 MUX2X1_14/a_30_54# MUX2X1_14/a_2_10# INVX2_12/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4454 MUX2X1_14/a_17_10# NOR2X1_1/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4455 vdd OAI21X1_1/Y MUX2X1_14/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4456 MUX2X1_14/a_30_10# OAI21X1_1/Y INVX2_12/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4457 gnd OAI21X1_1/Y MUX2X1_14/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4458 vdd INVX2_10/A MUX2X1_14/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4459 INVX2_12/A MUX2X1_14/a_2_10# MUX2X1_14/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4460 DFFSR_6/a_23_27# DFFSR_6/a_47_71# DFFSR_6/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4461 DFFSR_6/a_2_6# DFFSR_6/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4462 DFFSR_6/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4463 DFFSR_6/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4464 DFFSR_6/a_113_6# DFFSR_7/S DFFSR_6/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4465 DFFSR_6/a_10_61# DFFSR_6/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4466 DFFSR_6/a_113_6# DFFSR_6/a_47_4# DFFSR_6/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4467 vdd DFFSR_6/a_122_6# DFFSR_7/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4468 vdd DFFSR_7/S DFFSR_6/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4469 DFFSR_6/a_26_6# DFFSR_6/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4470 DFFSR_6/a_23_27# DFFSR_6/a_47_4# DFFSR_6/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4471 DFFSR_6/a_57_6# DFFSR_6/a_47_4# DFFSR_6/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4472 gnd DFFSR_6/a_10_61# DFFSR_6/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4473 DFFSR_6/a_105_6# DFFSR_6/a_47_4# DFFSR_6/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4474 vdd DFFSR_7/S DFFSR_6/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4475 gnd INVX2_0/A DFFSR_6/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4476 DFFSR_6/a_122_6# DFFSR_6/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4477 DFFSR_6/a_10_61# DFFSR_7/S DFFSR_6/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4478 gnd DFFSR_6/a_47_71# DFFSR_6/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4479 vdd DFFSR_6/R DFFSR_6/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4480 DFFSR_6/a_130_6# DFFSR_6/a_105_6# DFFSR_6/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4481 DFFSR_6/a_10_6# DFFSR_6/R DFFSR_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4482 vdd DFFSR_6/a_47_71# DFFSR_6/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4483 DFFSR_6/a_57_6# DFFSR_6/a_47_71# DFFSR_6/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4484 vdd INVX2_0/A DFFSR_6/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4485 vdd DFFSR_6/a_10_61# DFFSR_6/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4486 DFFSR_6/a_105_6# DFFSR_6/a_47_71# DFFSR_6/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4487 DFFSR_6/a_146_6# DFFSR_6/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4488 gnd DFFSR_6/a_122_6# DFFSR_7/D Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4489 DFFSR_6/a_113_6# DFFSR_6/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4490 DFFSR_6/a_113_6# DFFSR_6/a_47_71# DFFSR_6/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4491 gnd DFFSR_6/R DFFSR_6/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4492 gnd OAI22X1_6/A OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M4493 OAI22X1_0/a_2_6# INVX2_98/Y OAI22X1_0/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4494 OAI22X1_0/Y INVX2_91/Y OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4495 OAI22X1_0/Y INVX2_46/Y OAI22X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M4496 OAI22X1_0/a_28_54# INVX2_91/Y OAI22X1_0/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4497 OAI22X1_0/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4498 OAI22X1_0/a_2_6# INVX2_46/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4499 vdd INVX2_98/Y OAI22X1_0/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4500 NOR2X1_6/B OR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4501 NOR2X1_6/B OR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4502 INVX2_75/Y INVX2_75/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4503 INVX2_75/Y INVX2_75/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4504 INVX2_64/Y INVX2_64/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4505 INVX2_64/Y INVX2_64/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4506 INVX2_31/Y INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4507 INVX2_31/Y INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4508 INVX2_98/A INVX2_97/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4509 INVX2_98/A INVX2_97/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4510 INVX2_86/Y in_ans1[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4511 INVX2_86/Y in_ans1[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4512 INVX2_53/Y INVX2_53/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4513 INVX2_53/Y INVX2_53/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4514 INVX2_42/Y INVX2_42/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4515 INVX2_42/Y INVX2_42/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4516 gnd INVX2_19/A OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4517 vdd DFFSR_7/S INVX2_69/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4518 INVX2_69/A DFFSR_7/S OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4519 INVX2_69/A OAI21X1_5/A OAI21X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4520 OAI21X1_16/a_9_54# INVX2_19/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4521 OAI21X1_16/a_2_6# OAI21X1_5/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4522 gnd INVX2_8/Y XNOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4523 XNOR2X1_3/Y INVX2_8/Y XNOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4524 XNOR2X1_3/a_12_41# NOR2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4525 XNOR2X1_3/a_18_54# XNOR2X1_3/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4526 XNOR2X1_3/a_35_6# XNOR2X1_3/a_2_6# XNOR2X1_3/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4527 XNOR2X1_3/a_18_6# XNOR2X1_3/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4528 vdd INVX2_8/Y XNOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4529 vdd NOR2X1_1/Y XNOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4530 XNOR2X1_3/Y XNOR2X1_3/a_2_6# XNOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4531 XNOR2X1_3/a_35_54# INVX2_8/Y XNOR2X1_3/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4532 XNOR2X1_3/a_12_41# NOR2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4533 gnd NOR2X1_1/Y XNOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4534 AND2X2_3/a_2_6# NOR2X1_8/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4535 AND2X2_3/a_9_6# NOR2X1_8/B AND2X2_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M4536 AND2X2_3/Y AND2X2_3/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4537 AND2X2_3/Y AND2X2_3/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4538 vdd AND2X2_3/B AND2X2_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4539 gnd AND2X2_3/B AND2X2_3/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4540 NOR2X1_19/Y NOR2X1_19/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M4541 NOR2X1_19/Y NOR2X1_19/B NOR2X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M4542 NOR2X1_19/a_9_54# NOR2X1_19/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4543 gnd NOR2X1_19/B NOR2X1_19/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4544 gnd DFFSR_2/D MUX2X1_15/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4545 MUX2X1_15/a_17_50# DFFSR_2/D vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4546 INVX2_13/A OAI21X1_1/Y MUX2X1_15/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4547 MUX2X1_15/a_30_54# MUX2X1_15/a_2_10# INVX2_13/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4548 MUX2X1_15/a_17_10# DFFSR_2/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4549 vdd OAI21X1_1/Y MUX2X1_15/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4550 MUX2X1_15/a_30_10# OAI21X1_1/Y INVX2_13/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4551 gnd OAI21X1_1/Y MUX2X1_15/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4552 vdd DFFSR_2/D MUX2X1_15/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4553 INVX2_13/A MUX2X1_15/a_2_10# MUX2X1_15/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4554 DFFSR_7/a_23_27# DFFSR_7/a_47_71# DFFSR_7/a_2_6# vdd pfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4555 DFFSR_7/a_2_6# DFFSR_7/R vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4556 DFFSR_7/a_47_71# BUFX2_1/Y vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4557 DFFSR_7/a_47_71# BUFX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4558 DFFSR_7/a_113_6# DFFSR_7/S DFFSR_7/a_146_6# Gnd nfet w=20 l=2
+  ad=0.17n pd=82u as=80p ps=48u
M4559 DFFSR_7/a_10_61# DFFSR_7/a_23_27# vdd vdd pfet w=20 l=2
+  ad=0.17n pd=82u as=0 ps=0
M4560 DFFSR_7/a_113_6# DFFSR_7/a_47_4# DFFSR_7/a_105_6# vdd pfet w=10 l=2
+  ad=0.17n pd=82u as=59.999996p ps=32u
M4561 vdd DFFSR_7/a_122_6# INVX2_1/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4562 vdd DFFSR_7/S DFFSR_7/a_113_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4563 DFFSR_7/a_26_6# DFFSR_7/a_23_27# gnd Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0 ps=0
M4564 DFFSR_7/a_23_27# DFFSR_7/a_47_4# DFFSR_7/a_2_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4565 DFFSR_7/a_57_6# DFFSR_7/a_47_4# DFFSR_7/a_23_27# vdd pfet w=10 l=2
+  ad=0.11n pd=52u as=0 ps=0
M4566 gnd DFFSR_7/a_10_61# DFFSR_7/a_10_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4567 DFFSR_7/a_105_6# DFFSR_7/a_47_4# DFFSR_7/a_10_61# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0.17n ps=82u
M4568 vdd DFFSR_7/S DFFSR_7/a_10_61# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4569 gnd DFFSR_7/D DFFSR_7/a_57_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=59.999996p ps=32u
M4570 DFFSR_7/a_122_6# DFFSR_7/a_105_6# vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4571 DFFSR_7/a_10_61# DFFSR_7/S DFFSR_7/a_26_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4572 gnd DFFSR_7/a_47_71# DFFSR_7/a_47_4# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4573 vdd DFFSR_7/R DFFSR_7/a_122_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4574 DFFSR_7/a_130_6# DFFSR_7/a_105_6# DFFSR_7/a_122_6# Gnd nfet w=20 l=2
+  ad=80p pd=48u as=0.12n ps=52u
M4575 DFFSR_7/a_10_6# DFFSR_7/R DFFSR_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4576 vdd DFFSR_7/a_47_71# DFFSR_7/a_47_4# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4577 DFFSR_7/a_57_6# DFFSR_7/a_47_71# DFFSR_7/a_23_27# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4578 vdd DFFSR_7/D DFFSR_7/a_57_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4579 vdd DFFSR_7/a_10_61# DFFSR_7/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4580 DFFSR_7/a_105_6# DFFSR_7/a_47_71# DFFSR_7/a_10_61# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4581 DFFSR_7/a_146_6# DFFSR_7/a_122_6# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4582 gnd DFFSR_7/a_122_6# INVX2_1/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4583 DFFSR_7/a_113_6# DFFSR_7/a_122_6# vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4584 DFFSR_7/a_113_6# DFFSR_7/a_47_71# DFFSR_7/a_105_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4585 gnd DFFSR_7/R DFFSR_7/a_130_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4586 gnd OAI22X1_6/A OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M4587 OAI22X1_1/a_2_6# INVX2_98/Y OAI22X1_1/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4588 OAI22X1_1/Y INVX2_92/Y OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4589 OAI22X1_1/Y INVX2_45/Y OAI22X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M4590 OAI22X1_1/a_28_54# INVX2_92/Y OAI22X1_1/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4591 OAI22X1_1/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4592 OAI22X1_1/a_2_6# INVX2_45/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4593 vdd INVX2_98/Y OAI22X1_1/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4594 NOR2X1_1/B INVX2_10/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4595 NOR2X1_1/B INVX2_10/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4596 NOR2X1_7/B INVX2_21/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4597 NOR2X1_7/B INVX2_21/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4598 INVX2_65/Y INVX2_65/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4599 INVX2_65/Y INVX2_65/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4600 INVX2_76/Y INVX2_76/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4601 INVX2_76/Y INVX2_76/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4602 INVX2_98/Y INVX2_98/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4603 INVX2_98/Y INVX2_98/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4604 INVX2_32/Y INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4605 INVX2_32/Y INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4606 INVX2_87/Y in_ans1[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4607 INVX2_87/Y in_ans1[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4608 INVX2_43/Y INVX2_43/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4609 INVX2_43/Y INVX2_43/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4610 INVX2_54/Y INVX2_54/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4611 INVX2_54/Y INVX2_54/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4612 gnd OAI21X1_17/A OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4613 vdd AOI22X1_5/Y XOR2X1_3/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4614 XOR2X1_3/B AOI22X1_5/Y OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4615 XOR2X1_3/B OAI21X1_17/B OAI21X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4616 OAI21X1_17/a_9_54# OAI21X1_17/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4617 OAI21X1_17/a_2_6# OAI21X1_17/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4618 gnd INVX2_7/Y XNOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4619 MUX2X1_9/A INVX2_7/Y XNOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4620 XNOR2X1_4/a_12_41# INVX2_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4621 XNOR2X1_4/a_18_54# XNOR2X1_4/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4622 XNOR2X1_4/a_35_6# XNOR2X1_4/a_2_6# MUX2X1_9/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4623 XNOR2X1_4/a_18_6# XNOR2X1_4/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4624 vdd INVX2_7/Y XNOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4625 vdd INVX2_6/Y XNOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4626 MUX2X1_9/A XNOR2X1_4/a_2_6# XNOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4627 XNOR2X1_4/a_35_54# INVX2_7/Y MUX2X1_9/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4628 XNOR2X1_4/a_12_41# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4629 gnd INVX2_6/Y XNOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4630 AND2X2_4/a_2_6# INVX2_94/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4631 AND2X2_4/a_9_6# INVX2_94/Y AND2X2_4/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M4632 AND2X2_4/Y AND2X2_4/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4633 AND2X2_4/Y AND2X2_4/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4634 vdd AND2X2_4/B AND2X2_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4635 gnd AND2X2_4/B AND2X2_4/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4636 gnd XNOR2X1_1/Y MUX2X1_16/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4637 MUX2X1_16/a_17_50# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4638 INVX2_14/A OAI21X1_0/Y MUX2X1_16/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4639 MUX2X1_16/a_30_54# MUX2X1_16/a_2_10# INVX2_14/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4640 MUX2X1_16/a_17_10# INVX2_11/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4641 vdd OAI21X1_0/Y MUX2X1_16/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4642 MUX2X1_16/a_30_10# OAI21X1_0/Y INVX2_14/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4643 gnd OAI21X1_0/Y MUX2X1_16/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4644 vdd XNOR2X1_1/Y MUX2X1_16/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4645 INVX2_14/A MUX2X1_16/a_2_10# MUX2X1_16/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4646 OAI21X1_20/B XNOR2X1_68/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4647 NAND2X1_20/a_9_6# XNOR2X1_68/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4648 vdd XNOR2X1_67/Y OAI21X1_20/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4649 OAI21X1_20/B XNOR2X1_67/Y NAND2X1_20/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4650 gnd OAI22X1_6/A OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M4651 OAI22X1_2/a_2_6# INVX2_98/Y OAI22X1_2/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4652 OAI22X1_2/Y INVX2_93/Y OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4653 OAI22X1_2/Y INVX2_44/Y OAI22X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M4654 OAI22X1_2/a_28_54# INVX2_93/Y OAI22X1_2/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4655 OAI22X1_2/a_9_54# OAI22X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4656 OAI22X1_2/a_2_6# INVX2_44/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4657 vdd INVX2_98/Y OAI22X1_2/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4658 INVX2_11/Y INVX2_11/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4659 INVX2_11/Y INVX2_11/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4660 NOR2X1_8/B NOR2X1_9/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4661 NOR2X1_8/B NOR2X1_9/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4662 INVX2_33/Y INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4663 INVX2_33/Y INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4664 INVX2_44/Y INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4665 INVX2_44/Y INVX2_44/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4666 DFFSR_7/S INVX2_99/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4667 DFFSR_7/S INVX2_99/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4668 INVX2_77/Y INVX2_77/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4669 INVX2_77/Y INVX2_77/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4670 INVX2_66/Y NOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4671 INVX2_66/Y NOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4672 INVX2_88/Y in_ans1[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4673 INVX2_88/Y in_ans1[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4674 INVX2_55/Y INVX2_55/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4675 INVX2_55/Y INVX2_55/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4676 gnd OAI21X1_18/A OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4677 vdd AOI22X1_6/Y XOR2X1_5/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4678 XOR2X1_5/B AOI22X1_6/Y OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4679 XOR2X1_5/B OAI21X1_18/B OAI21X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4680 OAI21X1_18/a_9_54# OAI21X1_18/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4681 OAI21X1_18/a_2_6# OAI21X1_18/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4682 gnd INVX2_5/Y XNOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4683 MUX2X1_8/A INVX2_5/Y XNOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4684 XNOR2X1_5/a_12_41# NOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4685 XNOR2X1_5/a_18_54# XNOR2X1_5/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4686 XNOR2X1_5/a_35_6# XNOR2X1_5/a_2_6# MUX2X1_8/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4687 XNOR2X1_5/a_18_6# XNOR2X1_5/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4688 vdd INVX2_5/Y XNOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4689 vdd NOR2X1_2/Y XNOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4690 MUX2X1_8/A XNOR2X1_5/a_2_6# XNOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4691 XNOR2X1_5/a_35_54# INVX2_5/Y MUX2X1_8/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4692 XNOR2X1_5/a_12_41# NOR2X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4693 gnd NOR2X1_2/Y XNOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd OAI22X1_6/A 6.19641f
C1 XOR2X1_3/B vdd 2.16063f
C2 vdd INVX2_102/Y 15.225024f
C3 vdd INVX2_57/Y 3.1689f
C4 vdd INVX2_99/A 2.88576f
C5 vdd INVX2_33/A 3.15153f
C6 gnd INVX2_45/A 2.02239f
C7 OAI21X1_0/Y vdd 4.34079f
C8 vdd INVX2_1/A 2.93724f
C9 vdd INVX2_24/A 3.060451f
C10 vdd INVX2_44/A 3.036151f
C11 vdd OAI21X1_1/Y 4.85631f
C12 vdd INVX2_72/Y 6.76656f
C13 vdd OAI22X1_9/D 2.08188f
C14 vdd INVX2_0/A 2.41632f
C15 vdd INVX2_69/Y 2.35629f
C16 vdd OAI22X1_7/D 2.35431f
C17 vdd BUFX2_1/Y 2.23182f
C18 INVX2_40/A vdd 2.01492f
C19 vdd OAI21X1_17/B 2.16567f
C20 vdd INVX2_69/A 2.29761f
C21 vdd INVX2_39/Y 2.5524f
C22 vdd OR2X1_0/B 3.05892f
C23 INVX2_46/A vdd 4.80825f
C24 gnd INVX2_102/Y 2.820151f
C25 vdd INVX2_35/A 2.52711f
C26 vdd INVX2_101/Y 15.111534f
C27 vdd NAND2X1_4/Y 2.47662f
C28 vdd INVX2_32/A 5.17914f
C29 vdd INVX2_18/A 3.68361f
C30 vdd NOR2X1_1/B 2.06964f
C31 vdd INVX2_33/Y 2.00106f
C32 vdd INVX2_54/Y 2.33406f
C33 vdd NOR2X1_32/Y 2.46222f
C34 vdd MUX2X1_7/S 4.65012f
C35 vdd INVX2_25/A 3.851551f
C36 vdd INVX2_98/Y 10.527566f
C37 vdd INVX2_38/A 2.73933f
C38 INVX2_50/A vdd 2.19699f
C39 gnd vdd 5.832f
C40 NAND3X1_8/A vdd 2.05434f
C41 vdd INVX2_37/A 3.834361f
C42 gnd INVX2_101/Y 2.2644f
C43 vdd NOR2X1_8/B 3.0942f
C44 INVX4_0/Y vdd 24.475048f
C45 vdd INVX2_36/A 4.32135f
C46 vdd NAND2X1_4/A 2.65203f
C47 vdd INVX2_29/A 4.229551f
C48 vdd INVX2_27/A 4.39083f
C49 vdd INVX2_40/Y 2.88963f
C50 NOR2X1_9/A vdd 2.18097f
C51 vdd NOR2X1_9/B 3.43935f
C52 vdd AND2X2_2/B 2.20248f
C53 NAND2X1_3/A vdd 3.27141f
C54 vdd INVX2_23/A 3.97323f
C55 vdd INVX2_21/A 3.94245f
C56 DFFSR_4/D vdd 2.32002f
C57 vdd out_state[1] 3.23559f
C58 vdd INVX2_31/A 4.11417f
C59 vdd INVX2_68/A 2.06199f
C60 INVX2_67/Y vdd 2.57859f
C61 INVX2_47/A vdd 2.769751f
C62 vdd INVX2_28/A 4.131451f
C63 vdd DFFSR_7/S 13.340425f
C64 INVX4_0/Y gnd 4.347001f
C65 vdd INVX2_45/A 2.95218f
C66 vdd INVX2_62/Y 2.08143f
C67 vdd NOR2X1_8/Y 2.30589f
C68 vdd INVX2_30/A 3.89727f
C69 vdd MUX2X1_9/S 4.099861f
C70 vdd INVX2_67/A 2.42865f
C71 vdd INVX2_73/Y 3.07062f
C72 vdd NOR2X1_5/Y 4.19058f
C73 vdd NAND2X1_2/A 2.77155f
C74 vdd NOR2X1_7/A 3.2526f
C75 vdd AOI22X1_3/C 3.11229f
C76 INVX2_26/A vdd 3.79107f
C77 XNOR2X1_22/A 0 14.968951f **FLOATING
C78 OAI22X1_1/Y 0 11.977739f **FLOATING
C79 INVX2_98/Y 0 0.148068p **FLOATING
C80 OAI22X1_6/A 0 0.118382p **FLOATING
C81 OAI21X1_17/B 0 13.862841f **FLOATING
C82 NOR2X1_31/Y 0 13.083219f **FLOATING
C83 INVX2_53/A 0 15.999812f **FLOATING
C84 XNOR2X1_68/Y 0 11.39817f **FLOATING
C85 XNOR2X1_46/Y 0 14.893711f **FLOATING
C86 NOR2X1_33/B 0 17.934448f **FLOATING
C87 OAI21X1_20/B 0 9.094799f **FLOATING
C88 NOR2X1_31/B 0 10.61427f **FLOATING
C89 INVX2_23/A 0 42.24479f **FLOATING
C90 INVX2_45/A 0 57.23187f **FLOATING
C91 OAI21X1_20/A 0 11.216021f **FLOATING
C92 AOI22X1_5/Y 0 12.54492f **FLOATING
C93 INVX2_30/A 0 55.17112f **FLOATING
C94 NAND3X1_8/B 0 16.67448f **FLOATING
C95 NOR2X1_15/Y 0 10.85184f **FLOATING
C96 NOR2X1_16/Y 0 11.317762f **FLOATING
C97 INVX2_29/A 0 48.584812f **FLOATING
C98 INVX2_48/A 0 29.470844f **FLOATING
C99 NOR2X1_25/A 0 20.222607f **FLOATING
C100 XNOR2X1_90/Y 0 9.926489f **FLOATING
C101 INVX2_39/Y 0 40.89861f **FLOATING
C102 NOR2X1_28/Y 0 11.547961f **FLOATING
C103 NOR2X1_21/B 0 11.891069f **FLOATING
C104 NOR2X1_34/A 0 14.95809f **FLOATING
C105 NOR2X1_29/A 0 11.17275f **FLOATING
C106 INVX2_81/Y 0 8.77056f **FLOATING
C107 NOR2X1_17/Y 0 24.2412f **FLOATING
C108 NOR2X1_29/B 0 8.655809f **FLOATING
C109 NOR2X1_27/Y 0 14.083712f **FLOATING
C110 OAI22X1_6/Y 0 9.322202f **FLOATING
C111 INVX2_55/Y 0 35.814323f **FLOATING
C112 INVX2_55/A 0 20.409903f **FLOATING
C113 INVX2_54/Y 0 44.208298f **FLOATING
C114 NOR2X1_23/B 0 11.172091f **FLOATING
C115 NOR2X1_22/A 0 10.43025f **FLOATING
C116 NOR2X1_24/B 0 12.921929f **FLOATING
C117 NOR2X1_25/Y 0 10.468202f **FLOATING
C118 NOR2X1_32/Y 0 18.113367f **FLOATING
C119 OAI22X1_5/Y 0 10.744381f **FLOATING
C120 NOR2X1_26/B 0 10.336769f **FLOATING
C121 INVX2_102/Y 0 0.178615p **FLOATING
C122 NOR2X1_26/A 0 9.349709f **FLOATING
C123 INVX2_56/A 0 21.56202f **FLOATING
C124 NOR2X1_32/B 0 12.279869f **FLOATING
C125 INVX2_33/Y 0 20.0543f **FLOATING
C126 INVX2_67/A 0 37.152702f **FLOATING
C127 OAI22X1_15/Y 0 11.322959f **FLOATING
C128 INVX2_36/Y 0 10.867799f **FLOATING
C129 INVX2_35/Y 0 10.52682f **FLOATING
C130 OAI22X1_23/Y 0 9.38928f **FLOATING
C131 INVX2_37/Y 0 12.45234f **FLOATING
C132 INVX2_31/Y 0 8.7471f **FLOATING
C133 INVX2_26/Y 0 8.47284f **FLOATING
C134 INVX2_71/A 0 41.214153f **FLOATING
C135 OAI22X1_18/Y 0 11.472659f **FLOATING
C136 INVX2_69/A 0 49.689167f **FLOATING
C137 BUFX2_1/Y 0 37.194736f **FLOATING
C138 OAI22X1_19/Y 0 11.27028f **FLOATING
C139 OAI22X1_12/Y 0 10.425718f **FLOATING
C140 OAI22X1_9/D 0 36.410873f **FLOATING
C141 INVX2_19/A 0 24.98802f **FLOATING
C142 OAI22X1_14/Y 0 10.72404f **FLOATING
C143 DFFSR_7/D 0 22.292582f **FLOATING
C144 INVX2_68/A 0 38.181225f **FLOATING
C145 NOR2X1_10/B 0 13.67481f **FLOATING
C146 INVX2_72/Y 0 62.65148f **FLOATING
C147 INVX2_28/Y 0 9.5475f **FLOATING
C148 MUX2X1_0/A 0 9.210508f **FLOATING
C149 DFFSR_5/D 0 22.136488f **FLOATING
C150 OAI22X1_13/Y 0 10.5564f **FLOATING
C151 NAND2X1_9/Y 0 13.944839f **FLOATING
C152 NAND2X1_2/A 0 40.97021f **FLOATING
C153 OAI21X1_14/A 0 10.220401f **FLOATING
C154 NAND2X1_4/A 0 49.327106f **FLOATING
C155 AND2X2_3/B 0 24.712736f **FLOATING
C156 MUX2X1_0/Y 0 13.345591f **FLOATING
C157 NAND2X1_9/B 0 8.835211f **FLOATING
C158 OAI21X1_10/Y 0 10.010519f **FLOATING
C159 INVX2_5/A 0 14.6481f **FLOATING
C160 DFFSR_2/D 0 16.400818f **FLOATING
C161 NOR2X1_9/Y 0 16.020061f **FLOATING
C162 NOR2X1_7/Y 0 10.80276f **FLOATING
C163 OAI21X1_8/C 0 12.72825f **FLOATING
C164 MUX2X1_9/S 0 34.515953f **FLOATING
C165 NOR2X1_8/B 0 33.65237f **FLOATING
C166 AND2X2_4/B 0 11.595449f **FLOATING
C167 INVX2_6/Y 0 24.93933f **FLOATING
C168 INVX2_9/A 0 8.348701f **FLOATING
C169 OAI21X1_7/Y 0 10.353721f **FLOATING
C170 NOR2X1_6/Y 0 10.886701f **FLOATING
C171 INVX2_65/Y 0 9.660359f **FLOATING
C172 INVX2_11/Y 0 16.02399f **FLOATING
C173 INVX2_11/A 0 13.151159f **FLOATING
C174 OAI21X1_21/Y 0 11.0163f **FLOATING
C175 INVX2_61/A 0 8.45601f **FLOATING
C176 INVX2_92/Y 0 6.43386f **FLOATING
C177 XNOR2X1_71/A 0 13.279713f **FLOATING
C178 XNOR2X1_74/Y 0 16.36569f **FLOATING
C179 INVX2_60/A 0 28.84839f **FLOATING
C180 OAI22X1_0/Y 0 12.9198f **FLOATING
C181 INVX2_87/Y 0 7.889639f **FLOATING
C182 OAI22X1_28/Y 0 11.572379f **FLOATING
C183 INVX2_37/A 0 41.25858f **FLOATING
C184 INVX2_51/Y 0 26.102459f **FLOATING
C185 OAI22X1_29/Y 0 12.919801f **FLOATING
C186 INVX2_84/Y 0 6.71106f **FLOATING
C187 OAI22X1_25/Y 0 10.444499f **FLOATING
C188 INVX4_0/A 0 7.527059f **FLOATING
C189 INVX2_80/Y 0 8.447159f **FLOATING
C190 AND2X2_0/Y 0 10.185149f **FLOATING
C191 INVX2_36/A 0 46.810177f **FLOATING
C192 NOR2X1_20/B 0 11.48757f **FLOATING
C193 INVX2_50/Y 0 29.183388f **FLOATING
C194 NAND3X1_9/A 0 10.25703f **FLOATING
C195 INVX2_32/A 0 65.31166f **FLOATING
C196 XNOR2X1_55/Y 0 9.62391f **FLOATING
C197 INVX2_31/A 0 67.99399f **FLOATING
C198 XOR2X1_4/Y 0 18.043919f **FLOATING
C199 INVX2_58/A 0 8.7135f **FLOATING
C200 INVX2_51/A 0 31.218565f **FLOATING
C201 INVX2_83/Y 0 6.77766f **FLOATING
C202 OAI22X1_24/Y 0 11.431561f **FLOATING
C203 XNOR2X1_43/Y 0 9.74601f **FLOATING
C204 INVX2_28/A 0 52.446304f **FLOATING
C205 NOR2X1_5/Y 0 29.893263f **FLOATING
C206 NOR2X1_5/A 0 12.18066f **FLOATING
C207 INVX2_1/A 0 39.28991f **FLOATING
C208 MUX2X1_4/Y 0 12.83538f **FLOATING
C209 INVX2_3/Y 0 20.09262f **FLOATING
C210 INVX2_6/A 0 14.813641f **FLOATING
C211 INVX2_4/Y 0 20.05455f **FLOATING
C212 MUX2X1_7/S 0 27.995699f **FLOATING
C213 XOR2X1_1/Y 0 10.544401f **FLOATING
C214 XOR2X1_2/Y 0 13.15515f **FLOATING
C215 INVX2_0/A 0 45.668003f **FLOATING
C216 INVX2_25/A 0 50.15564f **FLOATING
C217 XOR2X1_5/Y 0 14.22492f **FLOATING
C218 OAI21X1_19/B 0 10.931221f **FLOATING
C219 AOI22X1_7/Y 0 25.738796f **FLOATING
C220 XNOR2X1_45/Y 0 9.625949f **FLOATING
C221 XNOR2X1_86/Y 0 9.97629f **FLOATING
C222 NOR2X1_30/B 0 9.698849f **FLOATING
C223 INVX2_41/Y 0 44.992603f **FLOATING
C224 OAI22X1_8/Y 0 11.640779f **FLOATING
C225 INVX2_7/A 0 14.579301f **FLOATING
C226 MUX2X1_9/A 0 9.283529f **FLOATING
C227 INVX2_8/Y 0 18.149488f **FLOATING
C228 INVX2_5/Y 0 19.78287f **FLOATING
C229 INVX2_40/Y 0 41.145782f **FLOATING
C230 INVX2_29/Y 0 8.51034f **FLOATING
C231 INVX2_32/Y 0 9.547502f **FLOATING
C232 OAI22X1_17/Y 0 12.58386f **FLOATING
C233 OAI21X1_18/B 0 18.201359f **FLOATING
C234 NOR2X1_22/Y 0 15.335098f **FLOATING
C235 INVX2_33/A 0 40.60916f **FLOATING
C236 INVX2_18/A 0 46.82435f **FLOATING
C237 XNOR2X1_58/Y 0 13.29765f **FLOATING
C238 XNOR2X1_33/Y 0 11.50089f **FLOATING
C239 INVX2_27/A 0 60.11155f **FLOATING
C240 OAI22X1_31/Y 0 11.06808f **FLOATING
C241 NOR2X1_15/B 0 8.02395f **FLOATING
C242 INVX2_38/A 0 40.62151f **FLOATING
C243 INVX2_47/Y 0 19.971748f **FLOATING
C244 INVX2_93/Y 0 11.35422f **FLOATING
C245 NOR2X1_15/A 0 10.06683f **FLOATING
C246 INVX2_35/A 0 34.711456f **FLOATING
C247 OAI22X1_8/D 0 25.852856f **FLOATING
C248 NOR2X1_34/Y 0 17.035757f **FLOATING
C249 NOR2X1_25/B 0 9.81813f **FLOATING
C250 NOR2X1_17/A 0 10.27479f **FLOATING
C251 INVX2_25/Y 0 8.435101f **FLOATING
C252 DFFSR_3/D 0 21.254217f **FLOATING
C253 INVX2_8/A 0 14.32794f **FLOATING
C254 INVX2_10/A 0 13.146481f **FLOATING
C255 INVX2_12/A 0 8.550659f **FLOATING
C256 NOR2X1_1/Y 0 18.487804f **FLOATING
C257 NOR2X1_1/B 0 24.801271f **FLOATING
C258 OAI21X1_1/Y 0 34.55178f **FLOATING
C259 NOR2X1_0/B 0 20.81941f **FLOATING
C260 INVX2_15/A 0 10.233541f **FLOATING
C261 INVX2_69/Y 0 28.306675f **FLOATING
C262 INVX2_30/Y 0 8.671741f **FLOATING
C263 NAND3X1_3/B 0 9.830009f **FLOATING
C264 NAND3X1_3/A 0 9.95043f **FLOATING
C265 INVX2_76/A 0 8.414099f **FLOATING
C266 INVX2_16/Y 0 10.988699f **FLOATING
C267 INVX2_17/A 0 10.68786f **FLOATING
C268 NAND3X1_5/B 0 8.839411f **FLOATING
C269 NAND3X1_5/A 0 12.51309f **FLOATING
C270 OAI22X1_7/Y 0 9.9711f **FLOATING
C271 INVX2_44/A 0 37.74428f **FLOATING
C272 INVX2_38/Y 0 8.123341f **FLOATING
C273 INVX2_24/A 0 30.718836f **FLOATING
C274 OAI22X1_27/Y 0 11.846519f **FLOATING
C275 INVX2_52/A 0 22.11516f **FLOATING
C276 INVX2_49/A 0 14.759431f **FLOATING
C277 INVX2_49/Y 0 35.409153f **FLOATING
C278 OAI22X1_30/Y 0 10.4445f **FLOATING
C279 INVX2_85/Y 0 6.43386f **FLOATING
C280 INVX2_68/Y 0 22.699879f **FLOATING
C281 INVX2_27/Y 0 9.90234f **FLOATING
C282 XNOR2X1_12/Y 0 8.86281f **FLOATING
C283 INVX2_75/A 0 9.16986f **FLOATING
C284 NOR2X1_0/Y 0 14.994122f **FLOATING
C285 in_clka 0 12.64659f **FLOATING
C286 INVX2_74/Y 0 11.31396f **FLOATING
C287 OAI22X1_7/D 0 32.862778f **FLOATING
C288 NAND2X1_4/Y 0 34.852486f **FLOATING
C289 INVX2_57/Y 0 50.47529f **FLOATING
C290 INVX2_71/Y 0 20.572956f **FLOATING
C291 INVX2_34/A 0 17.328537f **FLOATING
C292 INVX2_77/A 0 9.356939f **FLOATING
C293 INVX2_17/Y 0 15.009001f **FLOATING
C294 BUFX2_1/A 0 30.069662f **FLOATING
C295 INVX2_14/A 0 14.2485f **FLOATING
C296 INVX2_94/Y 0 10.730879f **FLOATING
C297 out_state[0] 0 18.717989f **FLOATING
C298 INVX2_95/Y 0 9.45084f **FLOATING
C299 out_state[1] 0 20.29586f **FLOATING
C300 INVX2_62/Y 0 24.31095f **FLOATING
C301 INVX2_64/Y 0 12.977221f **FLOATING
C302 AOI22X1_3/C 0 45.433186f **FLOATING
C303 DFFSR_7/S 0 0.207862p **FLOATING
C304 INVX2_99/A 0 37.152317f **FLOATING
C305 INVX2_23/Y 0 20.886597f **FLOATING
C306 AND2X2_2/B 0 26.932335f **FLOATING
C307 NOR2X1_8/Y 0 28.298098f **FLOATING
C308 INVX2_70/A 0 22.421217f **FLOATING
C309 INVX2_66/Y 0 7.793519f **FLOATING
C310 OR2X1_0/B 0 37.795704f **FLOATING
C311 OAI21X1_12/Y 0 10.00062f **FLOATING
C312 OAI21X1_21/C 0 9.83508f **FLOATING
C313 AOI21X1_3/B 0 18.740189f **FLOATING
C314 NOR2X1_36/Y 0 8.19918f **FLOATING
C315 out_valid 0 13.223671f **FLOATING
C316 INVX2_65/A 0 21.75648f **FLOATING
C317 NOR2X1_13/Y 0 12.724257f **FLOATING
C318 OAI21X1_6/B 0 11.95188f **FLOATING
C319 INVX2_98/A 0 7.89498f **FLOATING
C320 INVX2_82/Y 0 7.61376f **FLOATING
C321 INVX2_97/A 0 23.320587f **FLOATING
C322 NOR2X1_8/A 0 15.894392f **FLOATING
C323 NOR2X1_9/B 0 26.081009f **FLOATING
C324 INVX2_101/Y 0 0.163332p **FLOATING
C325 NAND3X1_2/Y 0 11.66805f **FLOATING
C326 INVX2_73/Y 0 22.228989f **FLOATING
C327 NOR2X1_6/A 0 21.951153f **FLOATING
C328 INVX2_21/A 0 28.772188f **FLOATING
C329 NOR2X1_7/A 0 49.115704f **FLOATING
C330 OAI21X1_8/Y 0 11.882641f **FLOATING
C331 INVX2_63/Y 0 16.555622f **FLOATING
C332 vdd 0 8.850143p **FLOATING
C333 XNOR2X1_5/a_2_6# 0 6.77121f **FLOATING
C334 XNOR2X1_5/a_12_41# 0 7.905991f **FLOATING
C335 OAI21X1_18/a_2_6# 0 2.78652f **FLOATING
C336 OAI21X1_18/A 0 6.67272f **FLOATING
C337 INVX2_88/Y 0 11.63142f **FLOATING
C338 OAI22X1_2/a_2_6# 0 4.25172f **FLOATING
C339 INVX2_44/Y 0 18.976952f **FLOATING
C340 INVX2_50/A 0 30.656425f **FLOATING
C341 XNOR2X1_1/Y 0 9.86901f **FLOATING
C342 MUX2X1_16/a_2_10# 0 6.0456f **FLOATING
C343 INVX2_42/Y 0 43.961185f **FLOATING
C344 INVX2_46/Y 0 7.519139f **FLOATING
C345 AND2X2_4/a_2_6# 0 6.03567f **FLOATING
C346 XNOR2X1_4/a_2_6# 0 6.77121f **FLOATING
C347 XNOR2X1_4/a_12_41# 0 7.905991f **FLOATING
C348 OAI21X1_17/a_2_6# 0 2.78652f **FLOATING
C349 NOR2X1_7/B 0 17.78502f **FLOATING
C350 OAI22X1_1/a_2_6# 0 4.25172f **FLOATING
C351 INVX2_42/A 0 14.01651f **FLOATING
C352 DFFSR_7/a_113_6# 0 11.4484f **FLOATING
C353 DFFSR_7/a_57_6# 0 4.37568f **FLOATING
C354 DFFSR_7/a_2_6# 0 11.1683f **FLOATING
C355 DFFSR_7/a_122_6# 0 7.77216f **FLOATING
C356 DFFSR_7/a_105_6# 0 6.46851f **FLOATING
C357 DFFSR_7/a_47_4# 0 10.7332f **FLOATING
C358 DFFSR_7/a_47_71# 0 11.4524f **FLOATING
C359 DFFSR_7/a_23_27# 0 6.98631f **FLOATING
C360 DFFSR_7/a_10_61# 0 14.156f **FLOATING
C361 DFFSR_7/R 0 8.388269f **FLOATING
C362 MUX2X1_15/a_2_10# 0 6.0456f **FLOATING
C363 NOR2X1_19/Y 0 11.19084f **FLOATING
C364 INVX2_52/Y 0 35.197582f **FLOATING
C365 AND2X2_3/Y 0 9.98703f **FLOATING
C366 AND2X2_3/a_2_6# 0 6.03567f **FLOATING
C367 XNOR2X1_3/a_2_6# 0 6.77121f **FLOATING
C368 XNOR2X1_3/a_12_41# 0 7.905991f **FLOATING
C369 OAI21X1_16/a_2_6# 0 2.78652f **FLOATING
C370 OAI21X1_5/A 0 16.612532f **FLOATING
C371 INVX2_86/Y 0 11.20926f **FLOATING
C372 OAI22X1_0/a_2_6# 0 4.25172f **FLOATING
C373 DFFSR_6/a_113_6# 0 11.4484f **FLOATING
C374 DFFSR_6/a_57_6# 0 4.37568f **FLOATING
C375 DFFSR_6/a_2_6# 0 11.1683f **FLOATING
C376 DFFSR_6/a_122_6# 0 7.77216f **FLOATING
C377 DFFSR_6/a_105_6# 0 6.46851f **FLOATING
C378 DFFSR_6/a_47_4# 0 10.7332f **FLOATING
C379 DFFSR_6/a_47_71# 0 11.4524f **FLOATING
C380 DFFSR_6/a_23_27# 0 6.98631f **FLOATING
C381 DFFSR_6/a_10_61# 0 14.156f **FLOATING
C382 DFFSR_6/R 0 8.388269f **FLOATING
C383 MUX2X1_14/a_2_10# 0 6.0456f **FLOATING
C384 NOR2X1_29/Y 0 14.386316f **FLOATING
C385 AND2X2_2/Y 0 7.55139f **FLOATING
C386 AND2X2_2/a_2_6# 0 6.03567f **FLOATING
C387 OAI21X1_0/Y 0 31.986498f **FLOATING
C388 XNOR2X1_2/a_2_6# 0 6.77121f **FLOATING
C389 XNOR2X1_2/a_12_41# 0 7.905991f **FLOATING
C390 OAI21X1_15/a_2_6# 0 2.78652f **FLOATING
C391 AOI21X1_2/B 0 13.027141f **FLOATING
C392 DFFSR_5/a_113_6# 0 11.4484f **FLOATING
C393 DFFSR_5/a_57_6# 0 4.37568f **FLOATING
C394 DFFSR_5/a_2_6# 0 11.1683f **FLOATING
C395 DFFSR_5/a_122_6# 0 7.77216f **FLOATING
C396 DFFSR_5/a_105_6# 0 6.46851f **FLOATING
C397 DFFSR_5/a_47_4# 0 10.7332f **FLOATING
C398 DFFSR_5/a_47_71# 0 11.4524f **FLOATING
C399 DFFSR_5/a_23_27# 0 6.98631f **FLOATING
C400 DFFSR_5/a_10_61# 0 14.156f **FLOATING
C401 DFFSR_5/R 0 8.388269f **FLOATING
C402 XNOR2X1_2/Y 0 9.86901f **FLOATING
C403 MUX2X1_13/a_2_10# 0 6.0456f **FLOATING
C404 NOR2X1_28/B 0 9.69885f **FLOATING
C405 OR2X1_0/A 0 16.78611f **FLOATING
C406 AND2X2_1/a_2_6# 0 6.03567f **FLOATING
C407 BUFX2_0/Y 0 15.572491f **FLOATING
C408 XNOR2X1_1/a_2_6# 0 6.77121f **FLOATING
C409 XNOR2X1_1/a_12_41# 0 7.905991f **FLOATING
C410 AOI21X1_2/Y 0 10.64757f **FLOATING
C411 OAI21X1_14/a_2_6# 0 2.78652f **FLOATING
C412 DFFSR_4/D 0 24.314968f **FLOATING
C413 DFFSR_4/a_113_6# 0 11.4484f **FLOATING
C414 DFFSR_4/a_57_6# 0 4.37568f **FLOATING
C415 DFFSR_4/a_2_6# 0 11.1683f **FLOATING
C416 DFFSR_4/a_122_6# 0 7.77216f **FLOATING
C417 DFFSR_4/a_105_6# 0 6.46851f **FLOATING
C418 DFFSR_4/a_47_4# 0 10.7332f **FLOATING
C419 DFFSR_4/a_47_71# 0 11.4524f **FLOATING
C420 DFFSR_4/a_23_27# 0 6.98631f **FLOATING
C421 DFFSR_4/a_10_61# 0 14.156f **FLOATING
C422 DFFSR_4/R 0 8.388269f **FLOATING
C423 XNOR2X1_3/Y 0 9.86901f **FLOATING
C424 MUX2X1_12/a_2_10# 0 6.0456f **FLOATING
C425 NOR2X1_27/A 0 8.13114f **FLOATING
C426 NOR2X1_16/B 0 9.11337f **FLOATING
C427 AND2X2_0/a_2_6# 0 6.03567f **FLOATING
C428 NOR2X1_0/A 0 15.830972f **FLOATING
C429 XNOR2X1_0/a_2_6# 0 6.77121f **FLOATING
C430 XNOR2X1_0/a_12_41# 0 7.905991f **FLOATING
C431 NOR2X1_9/A 0 35.40828f **FLOATING
C432 OAI21X1_13/a_2_6# 0 2.78652f **FLOATING
C433 out_Anum[2] 0 4.33032f **FLOATING
C434 in_restart 0 3.64296f **FLOATING
C435 NOR2X1_24/A 0 10.47909f **FLOATING
C436 DFFSR_3/a_113_6# 0 11.4484f **FLOATING
C437 DFFSR_3/a_57_6# 0 4.37568f **FLOATING
C438 DFFSR_3/a_2_6# 0 11.1683f **FLOATING
C439 DFFSR_3/a_122_6# 0 7.77216f **FLOATING
C440 DFFSR_3/a_105_6# 0 6.46851f **FLOATING
C441 DFFSR_3/a_47_4# 0 10.7332f **FLOATING
C442 DFFSR_3/a_47_71# 0 11.4524f **FLOATING
C443 DFFSR_3/a_23_27# 0 6.98631f **FLOATING
C444 DFFSR_3/a_10_61# 0 14.156f **FLOATING
C445 DFFSR_3/R 0 8.388269f **FLOATING
C446 MUX2X1_11/a_2_10# 0 6.0456f **FLOATING
C447 NOR2X1_37/Y 0 13.1292f **FLOATING
C448 OAI21X1_12/a_2_6# 0 2.78652f **FLOATING
C449 DFFSR_2/a_113_6# 0 11.4484f **FLOATING
C450 DFFSR_2/a_57_6# 0 4.37568f **FLOATING
C451 DFFSR_2/a_2_6# 0 11.1683f **FLOATING
C452 DFFSR_2/a_122_6# 0 7.77216f **FLOATING
C453 DFFSR_2/a_105_6# 0 6.46851f **FLOATING
C454 DFFSR_2/a_47_4# 0 10.7332f **FLOATING
C455 DFFSR_2/a_47_71# 0 11.4524f **FLOATING
C456 DFFSR_2/a_23_27# 0 6.98631f **FLOATING
C457 DFFSR_2/a_10_61# 0 14.156f **FLOATING
C458 DFFSR_2/R 0 8.388269f **FLOATING
C459 MUX2X1_10/a_2_10# 0 6.0456f **FLOATING
C460 NOR2X1_14/Y 0 18.586798f **FLOATING
C461 OAI21X1_22/a_2_6# 0 2.78652f **FLOATING
C462 OAI21X1_11/a_2_6# 0 2.78652f **FLOATING
C463 DFFSR_1/a_113_6# 0 11.4484f **FLOATING
C464 DFFSR_1/a_57_6# 0 4.37568f **FLOATING
C465 DFFSR_1/a_2_6# 0 11.1683f **FLOATING
C466 DFFSR_1/a_122_6# 0 7.77216f **FLOATING
C467 DFFSR_1/a_105_6# 0 6.46851f **FLOATING
C468 DFFSR_1/a_47_4# 0 10.7332f **FLOATING
C469 DFFSR_1/a_47_71# 0 11.4524f **FLOATING
C470 DFFSR_1/a_23_27# 0 6.98631f **FLOATING
C471 DFFSR_1/a_10_61# 0 14.156f **FLOATING
C472 DFFSR_1/R 0 8.388269f **FLOATING
C473 OAI21X1_10/a_2_6# 0 2.78652f **FLOATING
C474 OAI21X1_21/a_2_6# 0 2.78652f **FLOATING
C475 in_loadtest 0 8.22144f **FLOATING
C476 INVX2_91/Y 0 10.36494f **FLOATING
C477 DFFSR_0/a_113_6# 0 11.4484f **FLOATING
C478 DFFSR_0/a_57_6# 0 4.37568f **FLOATING
C479 DFFSR_0/a_2_6# 0 11.1683f **FLOATING
C480 DFFSR_0/a_122_6# 0 7.77216f **FLOATING
C481 DFFSR_0/a_105_6# 0 6.46851f **FLOATING
C482 DFFSR_0/a_47_4# 0 10.7332f **FLOATING
C483 DFFSR_0/a_47_71# 0 11.4524f **FLOATING
C484 DFFSR_0/a_23_27# 0 6.98631f **FLOATING
C485 DFFSR_0/a_10_61# 0 14.156f **FLOATING
C486 DFFSR_0/R 0 8.388269f **FLOATING
C487 NOR2X1_23/Y 0 9.872161f **FLOATING
C488 NOR2X1_23/A 0 8.13114f **FLOATING
C489 OAI21X1_20/a_2_6# 0 2.78652f **FLOATING
C490 AOI22X1_8/Y 0 12.124681f **FLOATING
C491 INVX2_90/Y 0 9.97881f **FLOATING
C492 NAND2X1_3/A 0 44.947453f **FLOATING
C493 NOR2X1_22/B 0 9.11337f **FLOATING
C494 NOR2X1_33/Y 0 13.179229f **FLOATING
C495 NOR2X1_11/Y 0 19.217278f **FLOATING
C496 OAI22X1_19/a_2_6# 0 4.25172f **FLOATING
C497 XNOR2X1_69/Y 0 11.30847f **FLOATING
C498 NAND2X1_9/A 0 7.445039f **FLOATING
C499 NOR2X1_32/A 0 8.22831f **FLOATING
C500 NOR2X1_21/A 0 8.22831f **FLOATING
C501 XNOR2X1_82/Y 0 10.827869f **FLOATING
C502 OAI22X1_29/a_2_6# 0 4.25172f **FLOATING
C503 OAI22X1_18/a_2_6# 0 4.25172f **FLOATING
C504 OAI22X1_28/a_2_6# 0 4.25172f **FLOATING
C505 OAI22X1_17/a_2_6# 0 4.25172f **FLOATING
C506 NOR2X1_30/Y 0 9.55038f **FLOATING
C507 XNOR2X1_67/Y 0 8.59941f **FLOATING
C508 OAI21X1_7/B 0 10.161541f **FLOATING
C509 OAI22X1_27/a_2_6# 0 4.25172f **FLOATING
C510 OAI22X1_16/a_2_6# 0 4.25172f **FLOATING
C511 XNOR2X1_89/Y 0 10.86459f **FLOATING
C512 NOR2X1_11/A 0 12.26829f **FLOATING
C513 XNOR2X1_19/a_2_6# 0 6.77121f **FLOATING
C514 XNOR2X1_19/a_12_41# 0 7.905991f **FLOATING
C515 OAI21X1_7/C 0 6.87006f **FLOATING
C516 INVX2_16/A 0 13.43634f **FLOATING
C517 OAI22X1_26/a_2_6# 0 4.25172f **FLOATING
C518 OAI22X1_15/a_2_6# 0 4.25172f **FLOATING
C519 XNOR2X1_29/a_2_6# 0 6.77121f **FLOATING
C520 XNOR2X1_29/a_12_41# 0 7.905991f **FLOATING
C521 NOR2X1_11/B 0 8.34555f **FLOATING
C522 XNOR2X1_18/a_2_6# 0 6.77121f **FLOATING
C523 XNOR2X1_18/a_12_41# 0 7.905991f **FLOATING
C524 gnd 0 2.140928p **FLOATING
C525 OAI22X1_25/a_2_6# 0 4.25172f **FLOATING
C526 OAI22X1_14/a_2_6# 0 4.25172f **FLOATING
C527 INVX2_43/A 0 20.1267f **FLOATING
C528 XNOR2X1_56/Y 0 9.39009f **FLOATING
C529 XNOR2X1_28/a_2_6# 0 6.77121f **FLOATING
C530 XNOR2X1_28/a_12_41# 0 7.905991f **FLOATING
C531 XNOR2X1_39/a_2_6# 0 6.77121f **FLOATING
C532 XNOR2X1_39/a_12_41# 0 7.905991f **FLOATING
C533 XNOR2X1_17/a_2_6# 0 6.77121f **FLOATING
C534 XNOR2X1_17/a_12_41# 0 7.905991f **FLOATING
C535 DFFNEGX1_9/a_66_6# 0 6.40992f **FLOATING
C536 DFFNEGX1_9/a_23_6# 0 6.85692f **FLOATING
C537 DFFNEGX1_9/a_34_4# 0 4.93023f **FLOATING
C538 DFFNEGX1_9/a_2_6# 0 9.33504f **FLOATING
C539 OAI22X1_21/Y 0 14.33352f **FLOATING
C540 OAI22X1_24/a_2_6# 0 4.25172f **FLOATING
C541 OAI22X1_13/a_2_6# 0 4.25172f **FLOATING
C542 NOR2X1_6/B 0 5.88042f **FLOATING
C543 XNOR2X1_49/a_2_6# 0 6.77121f **FLOATING
C544 XNOR2X1_49/a_12_41# 0 7.905991f **FLOATING
C545 NOR2X1_17/B 0 8.02395f **FLOATING
C546 XNOR2X1_27/a_2_6# 0 6.77121f **FLOATING
C547 XNOR2X1_27/a_12_41# 0 7.905991f **FLOATING
C548 NOR2X1_20/A 0 8.13114f **FLOATING
C549 XNOR2X1_38/a_2_6# 0 6.77121f **FLOATING
C550 XNOR2X1_38/a_12_41# 0 7.905991f **FLOATING
C551 XNOR2X1_16/a_2_6# 0 6.77121f **FLOATING
C552 XNOR2X1_16/a_12_41# 0 7.905991f **FLOATING
C553 INVX2_9/Y 0 19.40892f **FLOATING
C554 DFFNEGX1_8/a_66_6# 0 6.40992f **FLOATING
C555 DFFNEGX1_8/a_23_6# 0 6.85692f **FLOATING
C556 DFFNEGX1_8/a_34_4# 0 4.93023f **FLOATING
C557 DFFNEGX1_8/a_2_6# 0 9.33504f **FLOATING
C558 OAI22X1_23/a_2_6# 0 4.25172f **FLOATING
C559 OAI22X1_12/a_2_6# 0 4.25172f **FLOATING
C560 XNOR2X1_48/a_2_6# 0 6.77121f **FLOATING
C561 XNOR2X1_48/a_12_41# 0 7.905991f **FLOATING
C562 NOR2X1_27/B 0 11.040872f **FLOATING
C563 XNOR2X1_59/a_2_6# 0 6.77121f **FLOATING
C564 XNOR2X1_59/a_12_41# 0 7.905991f **FLOATING
C565 XNOR2X1_37/a_2_6# 0 6.77121f **FLOATING
C566 XNOR2X1_37/a_12_41# 0 7.905991f **FLOATING
C567 NOR2X1_16/A 0 11.610721f **FLOATING
C568 XNOR2X1_26/a_2_6# 0 6.77121f **FLOATING
C569 XNOR2X1_26/a_12_41# 0 7.905991f **FLOATING
C570 NOR2X1_10/A 0 8.22831f **FLOATING
C571 XNOR2X1_15/a_2_6# 0 6.77121f **FLOATING
C572 XNOR2X1_15/a_12_41# 0 7.905991f **FLOATING
C573 INVX2_7/Y 0 19.642529f **FLOATING
C574 DFFNEGX1_7/a_66_6# 0 6.40992f **FLOATING
C575 DFFNEGX1_7/a_23_6# 0 6.85692f **FLOATING
C576 DFFNEGX1_7/a_34_4# 0 4.93023f **FLOATING
C577 DFFNEGX1_7/a_2_6# 0 9.33504f **FLOATING
C578 OAI22X1_22/a_2_6# 0 4.25172f **FLOATING
C579 INVX2_18/Y 0 10.044181f **FLOATING
C580 OAI22X1_11/a_2_6# 0 4.25172f **FLOATING
C581 NOR2X1_30/A 0 11.796329f **FLOATING
C582 OAI21X1_9/a_2_6# 0 2.78652f **FLOATING
C583 XNOR2X1_47/a_2_6# 0 6.77121f **FLOATING
C584 XNOR2X1_47/a_12_41# 0 7.905991f **FLOATING
C585 XNOR2X1_25/a_2_6# 0 6.77121f **FLOATING
C586 XNOR2X1_25/a_12_41# 0 7.905991f **FLOATING
C587 NOR2X1_19/A 0 8.13114f **FLOATING
C588 XNOR2X1_36/a_2_6# 0 6.77121f **FLOATING
C589 XNOR2X1_36/a_12_41# 0 7.905991f **FLOATING
C590 XNOR2X1_69/a_2_6# 0 6.77121f **FLOATING
C591 XNOR2X1_69/a_12_41# 0 7.905991f **FLOATING
C592 XNOR2X1_58/a_2_6# 0 6.77121f **FLOATING
C593 XNOR2X1_58/a_12_41# 0 7.905991f **FLOATING
C594 INVX2_47/A 0 30.42234f **FLOATING
C595 XNOR2X1_14/a_2_6# 0 6.77121f **FLOATING
C596 XNOR2X1_14/a_12_41# 0 7.905991f **FLOATING
C597 OAI21X1_5/B 0 7.74018f **FLOATING
C598 DFFNEGX1_6/a_66_6# 0 6.40992f **FLOATING
C599 DFFNEGX1_6/a_23_6# 0 6.85692f **FLOATING
C600 DFFNEGX1_6/a_34_4# 0 4.93023f **FLOATING
C601 DFFNEGX1_6/a_2_6# 0 9.33504f **FLOATING
C602 OAI22X1_32/a_2_6# 0 4.25172f **FLOATING
C603 OAI22X1_10/a_2_6# 0 4.25172f **FLOATING
C604 INVX2_67/Y 0 21.051805f **FLOATING
C605 OAI22X1_21/a_2_6# 0 4.25172f **FLOATING
C606 OAI21X1_8/a_2_6# 0 2.78652f **FLOATING
C607 OR2X1_0/Y 0 10.094339f **FLOATING
C608 OR2X1_0/a_2_54# 0 6.27999f **FLOATING
C609 NOR2X1_3/Y 0 16.13946f **FLOATING
C610 XNOR2X1_79/a_2_6# 0 6.77121f **FLOATING
C611 XNOR2X1_79/a_12_41# 0 7.905991f **FLOATING
C612 XNOR2X1_68/a_2_6# 0 6.77121f **FLOATING
C613 XNOR2X1_68/a_12_41# 0 7.905991f **FLOATING
C614 NOR2X1_19/B 0 10.55547f **FLOATING
C615 XNOR2X1_35/a_2_6# 0 6.77121f **FLOATING
C616 XNOR2X1_35/a_12_41# 0 7.905991f **FLOATING
C617 XNOR2X1_24/a_2_6# 0 6.77121f **FLOATING
C618 XNOR2X1_24/a_12_41# 0 7.905991f **FLOATING
C619 XNOR2X1_46/a_2_6# 0 6.77121f **FLOATING
C620 XNOR2X1_46/a_12_41# 0 7.905991f **FLOATING
C621 XNOR2X1_57/Y 0 8.31795f **FLOATING
C622 XNOR2X1_57/a_2_6# 0 6.77121f **FLOATING
C623 XNOR2X1_57/a_12_41# 0 7.905991f **FLOATING
C624 XNOR2X1_13/Y 0 7.445039f **FLOATING
C625 XNOR2X1_13/a_2_6# 0 6.77121f **FLOATING
C626 XNOR2X1_13/a_12_41# 0 7.905991f **FLOATING
C627 INVX4_0/Y 0 0.243408p **FLOATING
C628 OAI21X1_4/B 0 9.49542f **FLOATING
C629 INVX2_14/Y 0 17.0475f **FLOATING
C630 DFFNEGX1_5/a_66_6# 0 6.40992f **FLOATING
C631 DFFNEGX1_5/a_23_6# 0 6.85692f **FLOATING
C632 DFFNEGX1_5/a_34_4# 0 4.93023f **FLOATING
C633 DFFNEGX1_5/a_2_6# 0 9.33504f **FLOATING
C634 OAI21X1_9/Y 0 13.604219f **FLOATING
C635 OAI22X1_31/a_2_6# 0 4.25172f **FLOATING
C636 OAI22X1_20/a_2_6# 0 4.25172f **FLOATING
C637 OAI21X1_7/a_2_6# 0 2.78652f **FLOATING
C638 INVX2_40/A 0 17.01579f **FLOATING
C639 XNOR2X1_89/a_2_6# 0 6.77121f **FLOATING
C640 XNOR2X1_89/a_12_41# 0 7.905991f **FLOATING
C641 XNOR2X1_78/a_2_6# 0 6.77121f **FLOATING
C642 XNOR2X1_78/a_12_41# 0 7.905991f **FLOATING
C643 XNOR2X1_67/a_2_6# 0 6.77121f **FLOATING
C644 XNOR2X1_67/a_12_41# 0 7.905991f **FLOATING
C645 XNOR2X1_45/a_2_6# 0 6.77121f **FLOATING
C646 XNOR2X1_45/a_12_41# 0 7.905991f **FLOATING
C647 XNOR2X1_34/Y 0 7.54221f **FLOATING
C648 XNOR2X1_34/a_2_6# 0 6.77121f **FLOATING
C649 XNOR2X1_34/a_12_41# 0 7.905991f **FLOATING
C650 XNOR2X1_56/a_2_6# 0 6.77121f **FLOATING
C651 XNOR2X1_56/a_12_41# 0 7.905991f **FLOATING
C652 XNOR2X1_23/a_2_6# 0 6.77121f **FLOATING
C653 XNOR2X1_23/a_12_41# 0 7.905991f **FLOATING
C654 XNOR2X1_12/a_2_6# 0 6.77121f **FLOATING
C655 XNOR2X1_12/a_12_41# 0 7.905991f **FLOATING
C656 DFFNEGX1_4/a_66_6# 0 6.40992f **FLOATING
C657 DFFNEGX1_4/a_23_6# 0 6.85692f **FLOATING
C658 DFFNEGX1_4/a_34_4# 0 4.93023f **FLOATING
C659 DFFNEGX1_4/a_2_6# 0 9.33504f **FLOATING
C660 OAI22X1_22/Y 0 11.942461f **FLOATING
C661 OAI22X1_30/a_2_6# 0 4.25172f **FLOATING
C662 XNOR2X1_85/Y 0 10.03113f **FLOATING
C663 OAI21X1_6/a_2_6# 0 2.78652f **FLOATING
C664 INVX2_70/Y 0 23.723059f **FLOATING
C665 XNOR2X1_66/a_2_6# 0 6.77121f **FLOATING
C666 XNOR2X1_66/a_12_41# 0 7.905991f **FLOATING
C667 XNOR2X1_88/a_2_6# 0 6.77121f **FLOATING
C668 XNOR2X1_88/a_12_41# 0 7.905991f **FLOATING
C669 XNOR2X1_44/Y 0 12.658831f **FLOATING
C670 XNOR2X1_44/a_2_6# 0 6.77121f **FLOATING
C671 XNOR2X1_44/a_12_41# 0 7.905991f **FLOATING
C672 NAND3X1_9/B 0 7.2603f **FLOATING
C673 XNOR2X1_77/a_2_6# 0 6.77121f **FLOATING
C674 XNOR2X1_77/a_12_41# 0 7.905991f **FLOATING
C675 XNOR2X1_33/a_2_6# 0 6.77121f **FLOATING
C676 XNOR2X1_33/a_12_41# 0 7.905991f **FLOATING
C677 out_Bnum[1] 0 4.99305f **FLOATING
C678 INVX2_58/Y 0 12.527189f **FLOATING
C679 XNOR2X1_22/a_2_6# 0 6.77121f **FLOATING
C680 XNOR2X1_22/a_12_41# 0 7.905991f **FLOATING
C681 XNOR2X1_55/a_2_6# 0 6.77121f **FLOATING
C682 XNOR2X1_55/a_12_41# 0 7.905991f **FLOATING
C683 XNOR2X1_11/a_2_6# 0 6.77121f **FLOATING
C684 XNOR2X1_11/a_12_41# 0 7.905991f **FLOATING
C685 AOI21X1_3/a_2_54# 0 4.3068f **FLOATING
C686 MUX2X1_9/a_2_10# 0 6.0456f **FLOATING
C687 DFFNEGX1_3/a_66_6# 0 6.40992f **FLOATING
C688 DFFNEGX1_3/a_23_6# 0 6.85692f **FLOATING
C689 DFFNEGX1_3/a_34_4# 0 4.93023f **FLOATING
C690 DFFNEGX1_3/a_2_6# 0 9.33504f **FLOATING
C691 OAI21X1_5/a_2_6# 0 2.78652f **FLOATING
C692 XNOR2X1_54/a_2_6# 0 6.77121f **FLOATING
C693 XNOR2X1_54/a_12_41# 0 7.905991f **FLOATING
C694 XNOR2X1_65/a_2_6# 0 6.77121f **FLOATING
C695 XNOR2X1_65/a_12_41# 0 7.905991f **FLOATING
C696 NOR2X1_34/B 0 8.34555f **FLOATING
C697 XNOR2X1_87/a_2_6# 0 6.77121f **FLOATING
C698 XNOR2X1_87/a_12_41# 0 7.905991f **FLOATING
C699 XNOR2X1_32/a_2_6# 0 6.77121f **FLOATING
C700 XNOR2X1_32/a_12_41# 0 7.905991f **FLOATING
C701 XNOR2X1_43/a_2_6# 0 6.77121f **FLOATING
C702 XNOR2X1_43/a_12_41# 0 7.905991f **FLOATING
C703 NOR2X1_31/A 0 8.22831f **FLOATING
C704 XNOR2X1_76/a_2_6# 0 6.77121f **FLOATING
C705 XNOR2X1_76/a_12_41# 0 7.905991f **FLOATING
C706 XNOR2X1_21/a_2_6# 0 6.77121f **FLOATING
C707 XNOR2X1_21/a_12_41# 0 7.905991f **FLOATING
C708 XNOR2X1_10/a_2_6# 0 6.77121f **FLOATING
C709 XNOR2X1_10/a_12_41# 0 7.905991f **FLOATING
C710 AOI21X1_2/a_2_54# 0 4.3068f **FLOATING
C711 INVX2_2/Y 0 16.200512f **FLOATING
C712 NOR2X1_18/Y 0 14.101199f **FLOATING
C713 NOR2X1_21/Y 0 10.920599f **FLOATING
C714 XNOR2X1_32/Y 0 11.64819f **FLOATING
C715 MUX2X1_8/Y 0 11.13726f **FLOATING
C716 MUX2X1_8/A 0 9.86901f **FLOATING
C717 MUX2X1_8/a_2_10# 0 6.0456f **FLOATING
C718 DFFNEGX1_2/a_66_6# 0 6.40992f **FLOATING
C719 DFFNEGX1_2/a_23_6# 0 6.85692f **FLOATING
C720 DFFNEGX1_2/a_34_4# 0 4.93023f **FLOATING
C721 DFFNEGX1_2/a_2_6# 0 9.33504f **FLOATING
C722 INVX2_75/Y 0 13.04382f **FLOATING
C723 OAI21X1_4/a_2_6# 0 2.78652f **FLOATING
C724 INVX2_26/A 0 58.64319f **FLOATING
C725 XNOR2X1_86/a_2_6# 0 6.77121f **FLOATING
C726 XNOR2X1_86/a_12_41# 0 7.905991f **FLOATING
C727 XNOR2X1_42/a_2_6# 0 6.77121f **FLOATING
C728 XNOR2X1_42/a_12_41# 0 7.905991f **FLOATING
C729 XNOR2X1_53/a_2_6# 0 6.77121f **FLOATING
C730 XNOR2X1_53/a_12_41# 0 7.905991f **FLOATING
C731 XNOR2X1_64/a_2_6# 0 6.77121f **FLOATING
C732 XNOR2X1_64/a_12_41# 0 7.905991f **FLOATING
C733 XNOR2X1_31/a_2_6# 0 6.77121f **FLOATING
C734 XNOR2X1_31/a_12_41# 0 7.905991f **FLOATING
C735 XNOR2X1_75/a_2_6# 0 6.77121f **FLOATING
C736 XNOR2X1_75/a_12_41# 0 7.905991f **FLOATING
C737 XNOR2X1_20/a_2_6# 0 6.77121f **FLOATING
C738 XNOR2X1_20/a_12_41# 0 7.905991f **FLOATING
C739 AOI21X1_1/Y 0 6.58671f **FLOATING
C740 AOI21X1_1/a_2_54# 0 4.3068f **FLOATING
C741 INVX2_1/Y 0 6.44484f **FLOATING
C742 BUFX2_1/a_2_6# 0 5.63946f **FLOATING
C743 INVX2_59/A 0 9.831841f **FLOATING
C744 DFFNEGX1_19/a_66_6# 0 6.40992f **FLOATING
C745 DFFNEGX1_19/a_23_6# 0 6.85692f **FLOATING
C746 DFFNEGX1_19/a_34_4# 0 4.93023f **FLOATING
C747 DFFNEGX1_19/a_2_6# 0 9.33504f **FLOATING
C748 MUX2X1_7/a_2_10# 0 6.0456f **FLOATING
C749 DFFNEGX1_1/a_66_6# 0 6.40992f **FLOATING
C750 DFFNEGX1_1/a_23_6# 0 6.85692f **FLOATING
C751 DFFNEGX1_1/a_34_4# 0 4.93023f **FLOATING
C752 DFFNEGX1_1/a_2_6# 0 9.33504f **FLOATING
C753 INVX2_76/Y 0 12.925019f **FLOATING
C754 INVX2_79/Y 0 7.70034f **FLOATING
C755 OAI21X1_3/a_2_6# 0 2.78652f **FLOATING
C756 XNOR2X1_52/a_2_6# 0 6.77121f **FLOATING
C757 XNOR2X1_52/a_12_41# 0 7.905991f **FLOATING
C758 XNOR2X1_63/a_2_6# 0 6.77121f **FLOATING
C759 XNOR2X1_63/a_12_41# 0 7.905991f **FLOATING
C760 XNOR2X1_85/a_2_6# 0 6.77121f **FLOATING
C761 XNOR2X1_85/a_12_41# 0 7.905991f **FLOATING
C762 INVX2_53/Y 0 6.60513f **FLOATING
C763 XNOR2X1_74/a_2_6# 0 6.77121f **FLOATING
C764 XNOR2X1_74/a_12_41# 0 7.905991f **FLOATING
C765 INVX2_60/Y 0 9.18888f **FLOATING
C766 XNOR2X1_41/a_2_6# 0 6.77121f **FLOATING
C767 XNOR2X1_41/a_12_41# 0 7.905991f **FLOATING
C768 NOR2X1_18/A 0 8.22831f **FLOATING
C769 XNOR2X1_30/a_2_6# 0 6.77121f **FLOATING
C770 XNOR2X1_30/a_12_41# 0 7.905991f **FLOATING
C771 AOI21X1_0/a_2_54# 0 4.3068f **FLOATING
C772 INVX2_73/A 0 16.809362f **FLOATING
C773 INVX2_74/A 0 8.134859f **FLOATING
C774 BUFX2_0/a_2_6# 0 5.63946f **FLOATING
C775 DFFNEGX1_29/a_66_6# 0 6.40992f **FLOATING
C776 DFFNEGX1_29/a_23_6# 0 6.85692f **FLOATING
C777 DFFNEGX1_29/a_34_4# 0 4.93023f **FLOATING
C778 DFFNEGX1_29/a_2_6# 0 9.33504f **FLOATING
C779 OAI22X1_2/Y 0 11.97774f **FLOATING
C780 DFFNEGX1_18/a_66_6# 0 6.40992f **FLOATING
C781 DFFNEGX1_18/a_23_6# 0 6.85692f **FLOATING
C782 DFFNEGX1_18/a_34_4# 0 4.93023f **FLOATING
C783 DFFNEGX1_18/a_2_6# 0 9.33504f **FLOATING
C784 OAI22X1_16/Y 0 11.54226f **FLOATING
C785 MUX2X1_6/a_2_10# 0 6.0456f **FLOATING
C786 XOR2X1_5/B 0 12.828481f **FLOATING
C787 XOR2X1_5/a_2_6# 0 8.278139f **FLOATING
C788 XOR2X1_5/a_13_43# 0 7.836241f **FLOATING
C789 DFFNEGX1_0/a_66_6# 0 6.40992f **FLOATING
C790 DFFNEGX1_0/a_23_6# 0 6.85692f **FLOATING
C791 DFFNEGX1_0/a_34_4# 0 4.93023f **FLOATING
C792 DFFNEGX1_0/a_2_6# 0 9.33504f **FLOATING
C793 INVX2_77/Y 0 13.04382f **FLOATING
C794 OAI21X1_2/a_2_6# 0 2.78652f **FLOATING
C795 NOR2X1_2/Y 0 16.775612f **FLOATING
C796 XNOR2X1_51/a_2_6# 0 6.77121f **FLOATING
C797 XNOR2X1_51/a_12_41# 0 7.905991f **FLOATING
C798 NOR2X1_28/A 0 8.22831f **FLOATING
C799 XNOR2X1_62/a_2_6# 0 6.77121f **FLOATING
C800 XNOR2X1_62/a_12_41# 0 7.905991f **FLOATING
C801 XNOR2X1_40/a_2_6# 0 6.77121f **FLOATING
C802 XNOR2X1_40/a_12_41# 0 7.905991f **FLOATING
C803 NAND3X1_8/A 0 14.69211f **FLOATING
C804 XNOR2X1_73/a_2_6# 0 6.77121f **FLOATING
C805 XNOR2X1_73/a_12_41# 0 7.905991f **FLOATING
C806 NOR2X1_33/A 0 8.13114f **FLOATING
C807 XNOR2X1_84/a_2_6# 0 6.77121f **FLOATING
C808 XNOR2X1_84/a_12_41# 0 7.905991f **FLOATING
C809 NOR2X1_18/B 0 9.55785f **FLOATING
C810 AOI22X1_6/Y 0 15.00741f **FLOATING
C811 DFFNEGX1_28/a_66_6# 0 6.40992f **FLOATING
C812 DFFNEGX1_28/a_23_6# 0 6.85692f **FLOATING
C813 DFFNEGX1_28/a_34_4# 0 4.93023f **FLOATING
C814 DFFNEGX1_28/a_2_6# 0 9.33504f **FLOATING
C815 DFFNEGX1_17/a_66_6# 0 6.40992f **FLOATING
C816 DFFNEGX1_17/a_23_6# 0 6.85692f **FLOATING
C817 DFFNEGX1_17/a_34_4# 0 4.93023f **FLOATING
C818 DFFNEGX1_17/a_2_6# 0 9.33504f **FLOATING
C819 DFFNEGX1_39/a_66_6# 0 6.40992f **FLOATING
C820 DFFNEGX1_39/a_23_6# 0 6.85692f **FLOATING
C821 DFFNEGX1_39/a_34_4# 0 4.93023f **FLOATING
C822 DFFNEGX1_39/a_2_6# 0 9.33504f **FLOATING
C823 XOR2X1_4/a_2_6# 0 8.278139f **FLOATING
C824 XOR2X1_4/a_13_43# 0 7.836241f **FLOATING
C825 MUX2X1_5/A 0 9.86901f **FLOATING
C826 MUX2X1_5/a_2_10# 0 6.0456f **FLOATING
C827 INVX2_78/Y 0 7.61376f **FLOATING
C828 OAI21X1_1/a_2_6# 0 2.78652f **FLOATING
C829 XNOR2X1_50/a_2_6# 0 6.77121f **FLOATING
C830 XNOR2X1_50/a_12_41# 0 7.905991f **FLOATING
C831 out_Anum[0] 0 4.99305f **FLOATING
C832 XNOR2X1_72/a_2_6# 0 6.77121f **FLOATING
C833 XNOR2X1_72/a_12_41# 0 7.905991f **FLOATING
C834 XNOR2X1_61/a_2_6# 0 6.77121f **FLOATING
C835 XNOR2X1_61/a_12_41# 0 7.905991f **FLOATING
C836 INVX2_56/Y 0 39.691685f **FLOATING
C837 XNOR2X1_83/a_2_6# 0 6.77121f **FLOATING
C838 XNOR2X1_83/a_12_41# 0 7.905991f **FLOATING
C839 DFFSR_0/D 0 11.79534f **FLOATING
C840 NOR2X1_26/Y 0 13.23396f **FLOATING
C841 DFFNEGX1_27/a_66_6# 0 6.40992f **FLOATING
C842 DFFNEGX1_27/a_23_6# 0 6.85692f **FLOATING
C843 DFFNEGX1_27/a_34_4# 0 4.93023f **FLOATING
C844 DFFNEGX1_27/a_2_6# 0 9.33504f **FLOATING
C845 OAI22X1_4/Y 0 11.97774f **FLOATING
C846 DFFNEGX1_38/a_66_6# 0 6.40992f **FLOATING
C847 DFFNEGX1_38/a_23_6# 0 6.85692f **FLOATING
C848 DFFNEGX1_38/a_34_4# 0 4.93023f **FLOATING
C849 DFFNEGX1_38/a_2_6# 0 9.33504f **FLOATING
C850 DFFNEGX1_16/a_66_6# 0 6.40992f **FLOATING
C851 DFFNEGX1_16/a_23_6# 0 6.85692f **FLOATING
C852 DFFNEGX1_16/a_34_4# 0 4.93023f **FLOATING
C853 DFFNEGX1_16/a_2_6# 0 9.33504f **FLOATING
C854 OAI22X1_11/Y 0 12.854639f **FLOATING
C855 MUX2X1_4/A 0 9.86901f **FLOATING
C856 MUX2X1_4/a_2_10# 0 6.0456f **FLOATING
C857 out_Bnum[0] 0 4.7571f **FLOATING
C858 XOR2X1_3/a_2_6# 0 8.278139f **FLOATING
C859 XOR2X1_3/a_13_43# 0 7.836241f **FLOATING
C860 OAI21X1_0/a_2_6# 0 2.78652f **FLOATING
C861 OAI21X1_0/C 0 11.202779f **FLOATING
C862 XNOR2X1_82/a_2_6# 0 6.77121f **FLOATING
C863 XNOR2X1_82/a_12_41# 0 7.905991f **FLOATING
C864 XNOR2X1_60/a_2_6# 0 6.77121f **FLOATING
C865 XNOR2X1_60/a_12_41# 0 7.905991f **FLOATING
C866 out_Anum[1] 0 4.99305f **FLOATING
C867 XNOR2X1_71/a_2_6# 0 6.77121f **FLOATING
C868 XNOR2X1_71/a_12_41# 0 7.905991f **FLOATING
C869 AOI22X1_8/a_2_54# 0 6.66f **FLOATING
C870 INVX2_46/A 0 55.755646f **FLOATING
C871 NOR2X1_10/Y 0 9.232679f **FLOATING
C872 DFFNEGX1_26/a_66_6# 0 6.40992f **FLOATING
C873 DFFNEGX1_26/a_23_6# 0 6.85692f **FLOATING
C874 DFFNEGX1_26/a_34_4# 0 4.93023f **FLOATING
C875 DFFNEGX1_26/a_2_6# 0 9.33504f **FLOATING
C876 DFFNEGX1_37/a_66_6# 0 6.40992f **FLOATING
C877 INVX2_54/A 0 8.28012f **FLOATING
C878 DFFNEGX1_37/a_23_6# 0 6.85692f **FLOATING
C879 DFFNEGX1_37/a_34_4# 0 4.93023f **FLOATING
C880 DFFNEGX1_37/a_2_6# 0 9.33504f **FLOATING
C881 OAI22X1_26/Y 0 11.58324f **FLOATING
C882 DFFNEGX1_15/a_66_6# 0 6.40992f **FLOATING
C883 DFFNEGX1_15/a_23_6# 0 6.85692f **FLOATING
C884 DFFNEGX1_15/a_34_4# 0 4.93023f **FLOATING
C885 DFFNEGX1_15/a_2_6# 0 9.33504f **FLOATING
C886 INVX2_4/A 0 14.235178f **FLOATING
C887 MUX2X1_3/a_2_10# 0 6.0456f **FLOATING
C888 XOR2X1_2/a_2_6# 0 8.278139f **FLOATING
C889 XOR2X1_2/a_13_43# 0 7.836241f **FLOATING
C890 XNOR2X1_81/Y 0 7.118729f **FLOATING
C891 XNOR2X1_81/a_2_6# 0 6.77121f **FLOATING
C892 XNOR2X1_81/a_12_41# 0 7.905991f **FLOATING
C893 XNOR2X1_70/Y 0 7.54221f **FLOATING
C894 XNOR2X1_70/a_2_6# 0 6.77121f **FLOATING
C895 XNOR2X1_70/a_12_41# 0 7.905991f **FLOATING
C896 AOI22X1_7/a_2_54# 0 6.66f **FLOATING
C897 NOR2X1_24/Y 0 12.29892f **FLOATING
C898 DFFNEGX1_25/a_66_6# 0 6.40992f **FLOATING
C899 DFFNEGX1_25/a_23_6# 0 6.85692f **FLOATING
C900 DFFNEGX1_25/a_34_4# 0 4.93023f **FLOATING
C901 DFFNEGX1_25/a_2_6# 0 9.33504f **FLOATING
C902 DFFNEGX1_36/a_66_6# 0 6.40992f **FLOATING
C903 DFFNEGX1_36/a_23_6# 0 6.85692f **FLOATING
C904 DFFNEGX1_36/a_34_4# 0 4.93023f **FLOATING
C905 DFFNEGX1_36/a_2_6# 0 9.33504f **FLOATING
C906 DFFNEGX1_14/a_66_6# 0 6.40992f **FLOATING
C907 DFFNEGX1_14/a_23_6# 0 6.85692f **FLOATING
C908 DFFNEGX1_14/a_34_4# 0 4.93023f **FLOATING
C909 DFFNEGX1_14/a_2_6# 0 9.33504f **FLOATING
C910 INVX2_3/A 0 8.27046f **FLOATING
C911 INVX2_0/Y 0 6.13938f **FLOATING
C912 MUX2X1_2/a_2_10# 0 6.0456f **FLOATING
C913 XOR2X1_1/a_2_6# 0 8.278139f **FLOATING
C914 XOR2X1_1/a_13_43# 0 7.836241f **FLOATING
C915 OAI22X1_9/a_2_6# 0 4.25172f **FLOATING
C916 XNOR2X1_80/a_2_6# 0 6.77121f **FLOATING
C917 XNOR2X1_80/a_12_41# 0 7.905991f **FLOATING
C918 AOI22X1_6/a_2_54# 0 6.66f **FLOATING
C919 OAI21X1_9/C 0 9.39765f **FLOATING
C920 DFFNEGX1_35/a_66_6# 0 6.40992f **FLOATING
C921 DFFNEGX1_35/a_23_6# 0 6.85692f **FLOATING
C922 DFFNEGX1_35/a_34_4# 0 4.93023f **FLOATING
C923 DFFNEGX1_35/a_2_6# 0 9.33504f **FLOATING
C924 DFFNEGX1_24/a_66_6# 0 6.40992f **FLOATING
C925 DFFNEGX1_24/a_23_6# 0 6.85692f **FLOATING
C926 DFFNEGX1_24/a_34_4# 0 4.93023f **FLOATING
C927 DFFNEGX1_24/a_2_6# 0 9.33504f **FLOATING
C928 DFFNEGX1_13/a_66_6# 0 6.40992f **FLOATING
C929 DFFNEGX1_13/a_23_6# 0 6.85692f **FLOATING
C930 DFFNEGX1_13/a_34_4# 0 4.93023f **FLOATING
C931 DFFNEGX1_13/a_2_6# 0 9.33504f **FLOATING
C932 INVX2_2/A 0 19.030499f **FLOATING
C933 MUX2X1_1/a_2_10# 0 6.0456f **FLOATING
C934 XOR2X1_0/a_2_6# 0 8.278139f **FLOATING
C935 XOR2X1_0/a_13_43# 0 7.836241f **FLOATING
C936 INVX2_39/A 0 8.28012f **FLOATING
C937 OAI22X1_8/a_2_6# 0 4.25172f **FLOATING
C938 INVX2_41/A 0 16.042831f **FLOATING
C939 XNOR2X1_90/a_2_6# 0 6.77121f **FLOATING
C940 XNOR2X1_90/a_12_41# 0 7.905991f **FLOATING
C941 OAI21X1_17/A 0 12.45024f **FLOATING
C942 AOI22X1_5/a_2_54# 0 6.66f **FLOATING
C943 NOR2X1_20/Y 0 14.342521f **FLOATING
C944 DFFNEGX1_34/a_66_6# 0 6.40992f **FLOATING
C945 DFFNEGX1_34/a_23_6# 0 6.85692f **FLOATING
C946 DFFNEGX1_34/a_34_4# 0 4.93023f **FLOATING
C947 DFFNEGX1_34/a_2_6# 0 9.33504f **FLOATING
C948 DFFNEGX1_12/a_66_6# 0 6.40992f **FLOATING
C949 DFFNEGX1_12/a_23_6# 0 6.85692f **FLOATING
C950 DFFNEGX1_12/a_34_4# 0 4.93023f **FLOATING
C951 DFFNEGX1_12/a_2_6# 0 9.33504f **FLOATING
C952 DFFNEGX1_23/a_66_6# 0 6.40992f **FLOATING
C953 DFFNEGX1_23/a_23_6# 0 6.85692f **FLOATING
C954 DFFNEGX1_23/a_34_4# 0 4.93023f **FLOATING
C955 DFFNEGX1_23/a_2_6# 0 9.33504f **FLOATING
C956 MUX2X1_0/a_2_10# 0 6.0456f **FLOATING
C957 OAI22X1_7/a_2_6# 0 4.25172f **FLOATING
C958 DFFSR_1/D 0 21.247442f **FLOATING
C959 AOI22X1_4/a_2_54# 0 6.66f **FLOATING
C960 XOR2X1_4/A 0 13.634731f **FLOATING
C961 XNOR2X1_31/Y 0 12.147209f **FLOATING
C962 DFFNEGX1_22/a_66_6# 0 6.40992f **FLOATING
C963 DFFNEGX1_22/a_23_6# 0 6.85692f **FLOATING
C964 DFFNEGX1_22/a_34_4# 0 4.93023f **FLOATING
C965 DFFNEGX1_22/a_2_6# 0 9.33504f **FLOATING
C966 OAI22X1_9/Y 0 11.28756f **FLOATING
C967 DFFNEGX1_33/a_66_6# 0 6.40992f **FLOATING
C968 DFFNEGX1_33/a_23_6# 0 6.85692f **FLOATING
C969 DFFNEGX1_33/a_34_4# 0 4.93023f **FLOATING
C970 DFFNEGX1_33/a_2_6# 0 9.33504f **FLOATING
C971 DFFNEGX1_11/a_66_6# 0 6.40992f **FLOATING
C972 DFFNEGX1_11/a_23_6# 0 6.85692f **FLOATING
C973 DFFNEGX1_11/a_34_4# 0 4.93023f **FLOATING
C974 DFFNEGX1_11/a_2_6# 0 9.33504f **FLOATING
C975 DFFNEGX1_44/a_66_6# 0 6.40992f **FLOATING
C976 DFFNEGX1_44/a_23_6# 0 6.85692f **FLOATING
C977 DFFNEGX1_44/a_34_4# 0 4.93023f **FLOATING
C978 DFFNEGX1_44/a_2_6# 0 9.33504f **FLOATING
C979 XNOR2X1_9/a_2_6# 0 6.77121f **FLOATING
C980 XNOR2X1_9/a_12_41# 0 7.905991f **FLOATING
C981 INVX2_64/A 0 11.83629f **FLOATING
C982 INVX2_48/Y 0 9.144481f **FLOATING
C983 out_Bnum[2] 0 4.33032f **FLOATING
C984 OAI22X1_6/a_2_6# 0 4.25172f **FLOATING
C985 XOR2X1_3/B 0 21.35634f **FLOATING
C986 AOI22X1_3/a_2_54# 0 6.66f **FLOATING
C987 INVX2_43/Y 0 19.79931f **FLOATING
C988 DFFNEGX1_21/a_66_6# 0 6.40992f **FLOATING
C989 DFFNEGX1_21/a_23_6# 0 6.85692f **FLOATING
C990 DFFNEGX1_21/a_34_4# 0 4.93023f **FLOATING
C991 DFFNEGX1_21/a_2_6# 0 9.33504f **FLOATING
C992 OAI22X1_10/Y 0 11.87892f **FLOATING
C993 DFFNEGX1_32/a_66_6# 0 6.40992f **FLOATING
C994 DFFNEGX1_32/a_23_6# 0 6.85692f **FLOATING
C995 DFFNEGX1_32/a_34_4# 0 4.93023f **FLOATING
C996 DFFNEGX1_32/a_2_6# 0 9.33504f **FLOATING
C997 DFFNEGX1_10/a_66_6# 0 6.40992f **FLOATING
C998 DFFNEGX1_10/a_23_6# 0 6.85692f **FLOATING
C999 DFFNEGX1_10/a_34_4# 0 4.93023f **FLOATING
C1000 DFFNEGX1_10/a_2_6# 0 9.33504f **FLOATING
C1001 OAI22X1_20/Y 0 13.38426f **FLOATING
C1002 DFFNEGX1_43/a_66_6# 0 6.40992f **FLOATING
C1003 DFFNEGX1_43/a_23_6# 0 6.85692f **FLOATING
C1004 DFFNEGX1_43/a_34_4# 0 4.93023f **FLOATING
C1005 DFFNEGX1_43/a_2_6# 0 9.33504f **FLOATING
C1006 MUX2X1_1/A 0 8.84631f **FLOATING
C1007 XNOR2X1_8/a_2_6# 0 6.77121f **FLOATING
C1008 XNOR2X1_8/a_12_41# 0 7.905991f **FLOATING
C1009 OAI22X1_5/a_2_6# 0 4.25172f **FLOATING
C1010 NOR2X1_37/B 0 10.002721f **FLOATING
C1011 AOI22X1_2/a_2_54# 0 6.66f **FLOATING
C1012 MUX2X1_19/a_2_10# 0 6.0456f **FLOATING
C1013 DFFNEGX1_31/a_66_6# 0 6.40992f **FLOATING
C1014 DFFNEGX1_31/a_23_6# 0 6.85692f **FLOATING
C1015 DFFNEGX1_31/a_34_4# 0 4.93023f **FLOATING
C1016 DFFNEGX1_31/a_2_6# 0 9.33504f **FLOATING
C1017 DFFNEGX1_20/a_66_6# 0 6.40992f **FLOATING
C1018 DFFNEGX1_20/a_23_6# 0 6.85692f **FLOATING
C1019 DFFNEGX1_20/a_34_4# 0 4.93023f **FLOATING
C1020 DFFNEGX1_20/a_2_6# 0 9.33504f **FLOATING
C1021 DFFNEGX1_42/a_66_6# 0 6.40992f **FLOATING
C1022 DFFNEGX1_42/a_23_6# 0 6.85692f **FLOATING
C1023 DFFNEGX1_42/a_34_4# 0 4.93023f **FLOATING
C1024 DFFNEGX1_42/a_2_6# 0 9.33504f **FLOATING
C1025 XNOR2X1_7/a_2_6# 0 6.77121f **FLOATING
C1026 XNOR2X1_7/a_12_41# 0 7.905991f **FLOATING
C1027 NOR2X1_35/Y 0 10.86438f **FLOATING
C1028 INVX2_57/A 0 8.235721f **FLOATING
C1029 INVX2_24/Y 0 14.54988f **FLOATING
C1030 OAI22X1_4/a_2_6# 0 4.25172f **FLOATING
C1031 AOI22X1_1/a_2_54# 0 6.66f **FLOATING
C1032 INVX2_15/Y 0 11.51274f **FLOATING
C1033 INVX2_13/A 0 11.942039f **FLOATING
C1034 MUX2X1_18/a_2_10# 0 6.0456f **FLOATING
C1035 DFFNEGX1_30/a_66_6# 0 6.40992f **FLOATING
C1036 DFFNEGX1_30/a_23_6# 0 6.85692f **FLOATING
C1037 DFFNEGX1_30/a_34_4# 0 4.93023f **FLOATING
C1038 DFFNEGX1_30/a_2_6# 0 9.33504f **FLOATING
C1039 DFFNEGX1_41/a_66_6# 0 6.40992f **FLOATING
C1040 DFFNEGX1_41/a_23_6# 0 6.85692f **FLOATING
C1041 DFFNEGX1_41/a_34_4# 0 4.93023f **FLOATING
C1042 DFFNEGX1_41/a_2_6# 0 9.33504f **FLOATING
C1043 AND2X2_4/Y 0 10.765351f **FLOATING
C1044 OAI22X1_3/Y 0 11.641981f **FLOATING
C1045 XNOR2X1_6/a_2_6# 0 6.77121f **FLOATING
C1046 XNOR2X1_6/a_12_41# 0 7.905991f **FLOATING
C1047 OAI21X1_19/a_2_6# 0 2.78652f **FLOATING
C1048 XOR2X1_5/A 0 12.858511f **FLOATING
C1049 OAI21X1_19/A 0 6.57834f **FLOATING
C1050 INVX2_89/Y 0 8.165999f **FLOATING
C1051 INVX2_45/Y 0 10.00722f **FLOATING
C1052 INVX2_34/Y 0 13.575361f **FLOATING
C1053 OAI22X1_3/a_2_6# 0 4.25172f **FLOATING
C1054 AOI22X1_0/a_2_54# 0 6.66f **FLOATING
C1055 XNOR2X1_0/Y 0 9.28353f **FLOATING
C1056 MUX2X1_17/a_2_10# 0 6.0456f **FLOATING
C1057 DFFNEGX1_40/a_66_6# 0 6.40992f **FLOATING
C1058 DFFNEGX1_40/a_23_6# 0 6.85692f **FLOATING
C1059 DFFNEGX1_40/a_34_4# 0 4.93023f **FLOATING
C1060 DFFNEGX1_40/a_2_6# 0 9.33504f **FLOATING
