* SPICE3 file created from hw5real.ext - technology: scmos

.option scale=0.15u

M1000 GND 17_14/DO 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1001 GND 17_14/a_26_538# 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1002 17_14/DATA 17_14/a_420_786# 17_14/DATA Gnd polyResistor w=20 l=128
+  ad=0.64n pd=0.104m as=1.618n ps=0.576m
M1003 17_14/DIB 17_14/DATA GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.378n ps=78u
M1004 17_14/a_62_902# 17_14/a_26_538# 17_14/a_62_82# Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0.624n ps=0.116m
M1005 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8n ps=0.28m
M1006 17_14/DI 17_14/DIB GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.378n ps=78u
M1007 Vdd 17_14/DO 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.648n pd=0.122m as=0.624n ps=0.116m
M1008 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.4n ps=0.284m
M1009 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.4n pd=0.284m as=3.6n ps=0.236m
M1010 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1011 Vdd 17_14/a_58_538# 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.648n pd=0.122m as=0.624n ps=0.116m
M1012 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8n pd=0.28m as=3.6n ps=0.236m
M1013 GND 17_14/a_26_538# 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.36n ps=72u
M1014 17_14/a_62_902# 17_14/a_58_538# 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.36n ps=72u
M1015 17_14/DIB 17_14/DATA Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.642n ps=0.122m
M1016 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.62n ps=0.44m
M1017 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M1018 17_14/a_62_82# 17_14/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.36n ps=72u
M1019 17_14/DI 17_14/DIB Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.642n ps=0.122m
M1020 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1021 17_14/a_62_82# 17_14/DO GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.378n ps=78u
M1022 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.708n pd=0.456m as=8.2n ps=0.282m
M1023 17_14/DATA 17_14/a_252_786# 17_14/DATA Gnd polyResistor w=20 l=130
+  ad=1.618n pd=0.576m as=0.6n ps=100u
M1024 Vdd 17_14/a_58_538# 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1025 17_14/a_62_82# 17_14/a_26_538# 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1026 GND 17_14/DATA 17_14/DIB Gnd nfet w=60 l=4
+  ad=0.378n pd=78u as=0.36n ps=72u
M1027 GND 17_14/DIB 17_14/DI Gnd nfet w=60 l=4
+  ad=0.378n pd=78u as=0.36n ps=72u
M1028 17_14/a_62_902# 17_14/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1029 17_14/a_62_902# 17_14/DO Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1030 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1031 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1032 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M1033 17_14/a_62_82# 17_14/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1034 17_14/a_62_82# 17_14/a_58_538# 17_14/a_62_902# Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.36n ps=72u
M1035 Vdd 17_14/DATA 17_14/DIB Vdd pfet w=104 l=4
+  ad=0.642n pd=0.122m as=0.624n ps=0.116m
M1036 Vdd 17_14/DIB 17_14/DI Vdd pfet w=104 l=4
+  ad=0.642n pd=0.122m as=0.624n ps=0.116m
M1037 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1038 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8n ps=0.28m
M1039 17_14/a_62_902# 17_14/a_26_538# 17_14/a_62_82# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1040 17_14/DIB 17_14/DATA GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1041 17_14/DI 17_14/DIB GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1042 17_14/a_62_902# 17_14/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.672n ps=0.128m
M1043 GND 17_14/DO 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.378n pd=78u as=0.72n ps=0.144m
M1044 GND 17_14/DO 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1045 17_14/a_58_538# 17_14/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0.36n ps=72u
M1046 17_14/a_62_902# 17_14/a_58_538# 17_14/a_62_82# Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.36n ps=72u
M1047 17_14/DI 17_14/DIB Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.648n ps=0.122m
M1048 Vdd 17_14/DO 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=1.248n ps=0.232m
M1049 17_14/DIB 17_14/DATA Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.648n ps=0.122m
M1050 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1051 17_14/DIB 17_14/DATA GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.78n ps=0.156m
M1052 17_14/DI 17_14/DIB GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1053 GND 17_14/DATA 17_14/DIB Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1054 17_14/a_58_538# 17_14/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0.624n ps=0.116m
M1055 Vdd 17_14/DO 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.672n pd=0.128m as=0.624n ps=0.116m
M1056 17_14/a_62_82# 17_14/a_26_538# 17_14/a_62_902# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.624n ps=0.116m
M1057 GND 17_14/DIB 17_14/DI Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1058 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1059 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8n pd=0.28m as=3.6n ps=0.236m
M1060 17_14/DIB 17_14/DATA Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=1.368n ps=0.256m
M1061 17_14/DI 17_14/DIB Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.672n ps=0.128m
M1062 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.4n ps=0.284m
M1063 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.4n pd=0.284m as=3.6n ps=0.236m
M1064 17_14/a_62_82# 17_14/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1065 GND 17_14/a_62_82# 17_14/DATA GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1066 GND 17_14/OEN 17_14/a_26_538# Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.72n ps=0.144m
M1067 17_14/a_62_82# 17_14/DO GND Gnd nfet w=60 l=4
+  ad=0.36n pd=72u as=0.384n ps=78u
M1068 Vdd 17_14/DATA 17_14/DIB Vdd pfet w=104 l=4
+  ad=0.648n pd=0.122m as=0.624n ps=0.116m
M1069 Vdd 17_14/DIB 17_14/DI Vdd pfet w=104 l=4
+  ad=0.648n pd=0.122m as=0.624n ps=0.116m
M1070 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1071 17_14/DATA 17_14/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M1072 Vdd 17_14/a_62_902# 17_14/DATA Vdd pfet w=200 l=6
+  ad=3.708n pd=0.456m as=8.2n ps=0.282m
M1073 GND 17_14/DATA 17_14/DIB Gnd nfet w=60 l=4
+  ad=0.384n pd=78u as=0.36n ps=72u
M1074 GND 17_14/DIB 17_14/DI Gnd nfet w=60 l=4
+  ad=0.648n pd=0.152m as=0.36n ps=72u
M1075 17_14/a_62_902# 17_14/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.648n ps=0.122m
M1076 Vdd 17_14/OEN 17_14/a_26_538# Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=1.248n ps=0.232m
M1077 17_14/a_62_902# 17_14/DO Vdd Vdd pfet w=104 l=4
+  ad=0.624n pd=0.116m as=0.648n ps=0.122m
M1078 17_14/a_62_82# 17_14/a_58_538# 17_14/a_62_902# Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0.36n ps=72u
M1079 Vdd 17_14/DATA 17_14/DIB Vdd pfet w=104 l=4
+  ad=0.672n pd=0.128m as=0.624n ps=0.116m
M1080 Vdd 17_14/DIB 17_14/DI Vdd pfet w=104 l=4
+  ad=1.28n pd=0.288m as=0.624n ps=0.116m
M1081 17_14/DATA 17_14/a_62_82# GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1082 GND 17_25/DO 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=1.994384u pd=0.210504 as=5.76n ps=1.152m
M1083 GND 17_25/a_26_538# 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1084 17_25/DATA 17_25/a_420_786# 17_25/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1085 17_25/DIB 17_25/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1086 17_25/a_62_902# 17_25/a_26_538# 17_25/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1087 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=2.256592u pd=0.25586 as=97.6n ps=3.376m
M1088 17_25/DI 17_25/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1089 Vdd 17_25/DO 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1090 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1091 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1092 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1093 Vdd 17_25/a_58_538# 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1094 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1095 GND 17_25/a_26_538# 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1096 17_25/a_62_902# 17_25/a_58_538# 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1097 17_25/DIB 17_25/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1098 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1099 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1100 17_25/a_62_82# 17_25/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1101 17_25/DI 17_25/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1102 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1103 17_25/a_62_82# 17_25/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1104 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1105 17_25/DATA 17_25/a_252_786# 17_25/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1106 Vdd 17_25/a_58_538# 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1107 17_25/a_62_82# 17_25/a_26_538# 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1108 GND 17_25/DATA 17_25/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1109 GND 17_25/DIB 17_25/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1110 17_25/a_62_902# 17_25/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1111 17_25/a_62_902# 17_25/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1113 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1114 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1115 17_25/a_62_82# 17_25/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1116 17_25/a_62_82# 17_25/a_58_538# 17_25/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1117 Vdd 17_25/DATA 17_25/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1118 Vdd 17_25/DIB 17_25/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1119 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1120 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1121 17_25/a_62_902# 17_25/a_26_538# 17_25/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1122 17_25/DIB 17_25/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1123 17_25/DI 17_25/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1124 17_25/a_62_902# 17_25/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1125 GND 17_25/DO 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1126 GND 17_25/DO 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1127 17_25/a_58_538# 17_25/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1128 17_25/a_62_902# 17_25/a_58_538# 17_25/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1129 17_25/DI 17_25/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 Vdd 17_25/DO 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1131 17_25/DIB 17_25/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1132 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1133 17_25/DIB 17_25/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1134 17_25/DI 17_25/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1135 GND 17_25/DATA 17_25/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1136 17_25/a_58_538# 17_25/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1137 Vdd 17_25/DO 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1138 17_25/a_62_82# 17_25/a_26_538# 17_25/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1139 GND 17_25/DIB 17_25/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1140 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1141 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1142 17_25/DIB 17_25/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1143 17_25/DI 17_25/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1144 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1145 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1146 17_25/a_62_82# 17_25/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1147 GND 17_25/a_62_82# 17_25/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1148 GND 17_25/OEN 17_25/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1149 17_25/a_62_82# 17_25/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1150 Vdd 17_25/DATA 17_25/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1151 Vdd 17_25/DIB 17_25/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1152 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1153 17_25/DATA 17_25/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1154 Vdd 17_25/a_62_902# 17_25/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1155 GND 17_25/DATA 17_25/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1156 GND 17_25/DIB 17_25/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1157 17_25/a_62_902# 17_25/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1158 Vdd 17_25/OEN 17_25/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1159 17_25/a_62_902# 17_25/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1160 17_25/a_62_82# 17_25/a_58_538# 17_25/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1161 Vdd 17_25/DATA 17_25/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1162 Vdd 17_25/DIB 17_25/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1163 17_25/DATA 17_25/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1164 GND 17_15/DO 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1165 GND 17_15/a_26_538# 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1166 17_15/DATA 17_15/a_420_786# 17_15/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1167 17_15/DIB 17_15/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1168 17_15/a_62_902# 17_15/a_26_538# 17_15/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1169 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1170 17_15/DI 17_15/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1171 Vdd 17_15/DO 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1172 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1173 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1174 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1175 Vdd 17_15/a_58_538# 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1176 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1177 GND 17_15/a_26_538# 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1178 17_15/a_62_902# 17_15/a_58_538# 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1179 17_15/DIB 17_15/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1180 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1181 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1182 17_15/a_62_82# 17_15/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1183 17_15/DI 17_15/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1184 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1185 17_15/a_62_82# 17_15/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1186 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1187 17_15/DATA 17_15/a_252_786# 17_15/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1188 Vdd 17_15/a_58_538# 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1189 17_15/a_62_82# 17_15/a_26_538# 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1190 GND 17_15/DATA 17_15/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1191 GND 17_15/DIB 17_15/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1192 17_15/a_62_902# 17_15/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1193 17_15/a_62_902# 17_15/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1194 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1195 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1196 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1197 17_15/a_62_82# 17_15/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1198 17_15/a_62_82# 17_15/a_58_538# 17_15/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1199 Vdd 17_15/DATA 17_15/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1200 Vdd 17_15/DIB 17_15/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1201 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1202 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1203 17_15/a_62_902# 17_15/a_26_538# 17_15/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1204 17_15/DIB 17_15/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1205 17_15/DI 17_15/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1206 17_15/a_62_902# 17_15/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1207 GND 17_15/DO 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1208 GND 17_15/DO 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1209 17_15/a_58_538# 17_15/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1210 17_15/a_62_902# 17_15/a_58_538# 17_15/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1211 17_15/DI 17_15/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1212 Vdd 17_15/DO 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1213 17_15/DIB 17_15/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1214 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1215 17_15/DIB 17_15/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1216 17_15/DI 17_15/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1217 GND 17_15/DATA 17_15/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1218 17_15/a_58_538# 17_15/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1219 Vdd 17_15/DO 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1220 17_15/a_62_82# 17_15/a_26_538# 17_15/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1221 GND 17_15/DIB 17_15/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1222 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1223 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1224 17_15/DIB 17_15/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1225 17_15/DI 17_15/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1226 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1227 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1228 17_15/a_62_82# 17_15/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1229 GND 17_15/a_62_82# 17_15/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1230 GND 17_15/OEN 17_15/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1231 17_15/a_62_82# 17_15/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1232 Vdd 17_15/DATA 17_15/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1233 Vdd 17_15/DIB 17_15/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1234 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1235 17_15/DATA 17_15/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1236 Vdd 17_15/a_62_902# 17_15/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1237 GND 17_15/DATA 17_15/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1238 GND 17_15/DIB 17_15/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1239 17_15/a_62_902# 17_15/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1240 Vdd 17_15/OEN 17_15/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1241 17_15/a_62_902# 17_15/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1242 17_15/a_62_82# 17_15/a_58_538# 17_15/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1243 Vdd 17_15/DATA 17_15/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1244 Vdd 17_15/DIB 17_15/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1245 17_15/DATA 17_15/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1246 GND 17_26/DO 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1247 GND 17_26/a_26_538# 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1248 17_26/DATA 17_26/a_420_786# 17_26/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1249 17_26/DIB 17_26/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1250 17_26/a_62_902# 17_26/a_26_538# 17_26/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1251 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1252 17_26/DI 17_26/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1253 Vdd 17_26/DO 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1254 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1255 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1256 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1257 Vdd 17_26/a_58_538# 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1258 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1259 GND 17_26/a_26_538# 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1260 17_26/a_62_902# 17_26/a_58_538# 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1261 17_26/DIB 17_26/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1262 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1263 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1264 17_26/a_62_82# 17_26/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1265 17_26/DI 17_26/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1266 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1267 17_26/a_62_82# 17_26/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1268 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1269 17_26/DATA 17_26/a_252_786# 17_26/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1270 Vdd 17_26/a_58_538# 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1271 17_26/a_62_82# 17_26/a_26_538# 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1272 GND 17_26/DATA 17_26/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1273 GND 17_26/DIB 17_26/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1274 17_26/a_62_902# 17_26/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1275 17_26/a_62_902# 17_26/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1276 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1277 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1278 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1279 17_26/a_62_82# 17_26/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1280 17_26/a_62_82# 17_26/a_58_538# 17_26/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1281 Vdd 17_26/DATA 17_26/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1282 Vdd 17_26/DIB 17_26/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1283 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1284 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1285 17_26/a_62_902# 17_26/a_26_538# 17_26/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1286 17_26/DIB 17_26/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1287 17_26/DI 17_26/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1288 17_26/a_62_902# 17_26/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1289 GND 17_26/DO 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1290 GND 17_26/DO 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1291 17_26/a_58_538# 17_26/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1292 17_26/a_62_902# 17_26/a_58_538# 17_26/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1293 17_26/DI 17_26/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1294 Vdd 17_26/DO 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1295 17_26/DIB 17_26/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1296 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1297 17_26/DIB 17_26/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1298 17_26/DI 17_26/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1299 GND 17_26/DATA 17_26/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1300 17_26/a_58_538# 17_26/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1301 Vdd 17_26/DO 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1302 17_26/a_62_82# 17_26/a_26_538# 17_26/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1303 GND 17_26/DIB 17_26/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1304 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1305 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1306 17_26/DIB 17_26/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1307 17_26/DI 17_26/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1308 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1309 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1310 17_26/a_62_82# 17_26/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1311 GND 17_26/a_62_82# 17_26/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1312 GND 17_26/OEN 17_26/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1313 17_26/a_62_82# 17_26/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1314 Vdd 17_26/DATA 17_26/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1315 Vdd 17_26/DIB 17_26/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1316 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1317 17_26/DATA 17_26/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1318 Vdd 17_26/a_62_902# 17_26/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1319 GND 17_26/DATA 17_26/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1320 GND 17_26/DIB 17_26/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1321 17_26/a_62_902# 17_26/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1322 Vdd 17_26/OEN 17_26/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1323 17_26/a_62_902# 17_26/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1324 17_26/a_62_82# 17_26/a_58_538# 17_26/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1325 Vdd 17_26/DATA 17_26/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1326 Vdd 17_26/DIB 17_26/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1327 17_26/DATA 17_26/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1328 GND 17_16/DO 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1329 GND 17_16/a_26_538# 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1330 17_16/DATA 17_16/a_420_786# 17_16/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1331 17_16/DIB 17_16/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1332 17_16/a_62_902# 17_16/a_26_538# 17_16/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1333 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1334 17_16/DI 17_16/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1335 Vdd 17_16/DO 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1336 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1337 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1338 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1339 Vdd 17_16/a_58_538# 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1340 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1341 GND 17_16/a_26_538# 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1342 17_16/a_62_902# 17_16/a_58_538# 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1343 17_16/DIB 17_16/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1344 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1345 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1346 17_16/a_62_82# 17_16/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1347 17_16/DI 17_16/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1348 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1349 17_16/a_62_82# 17_16/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1350 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1351 17_16/DATA 17_16/a_252_786# 17_16/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1352 Vdd 17_16/a_58_538# 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1353 17_16/a_62_82# 17_16/a_26_538# 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1354 GND 17_16/DATA 17_16/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1355 GND 17_16/DIB 17_16/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1356 17_16/a_62_902# 17_16/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1357 17_16/a_62_902# 17_16/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1358 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1359 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1360 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1361 17_16/a_62_82# 17_16/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1362 17_16/a_62_82# 17_16/a_58_538# 17_16/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1363 Vdd 17_16/DATA 17_16/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1364 Vdd 17_16/DIB 17_16/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1365 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1366 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1367 17_16/a_62_902# 17_16/a_26_538# 17_16/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1368 17_16/DIB 17_16/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1369 17_16/DI 17_16/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1370 17_16/a_62_902# 17_16/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1371 GND 17_16/DO 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1372 GND 17_16/DO 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1373 17_16/a_58_538# 17_16/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1374 17_16/a_62_902# 17_16/a_58_538# 17_16/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1375 17_16/DI 17_16/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1376 Vdd 17_16/DO 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1377 17_16/DIB 17_16/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1378 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1379 17_16/DIB 17_16/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1380 17_16/DI 17_16/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1381 GND 17_16/DATA 17_16/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1382 17_16/a_58_538# 17_16/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1383 Vdd 17_16/DO 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1384 17_16/a_62_82# 17_16/a_26_538# 17_16/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1385 GND 17_16/DIB 17_16/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1386 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1387 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1388 17_16/DIB 17_16/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1389 17_16/DI 17_16/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1390 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1391 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1392 17_16/a_62_82# 17_16/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1393 GND 17_16/a_62_82# 17_16/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1394 GND 17_16/OEN 17_16/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1395 17_16/a_62_82# 17_16/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1396 Vdd 17_16/DATA 17_16/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1397 Vdd 17_16/DIB 17_16/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1398 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1399 17_16/DATA 17_16/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1400 Vdd 17_16/a_62_902# 17_16/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1401 GND 17_16/DATA 17_16/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1402 GND 17_16/DIB 17_16/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1403 17_16/a_62_902# 17_16/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1404 Vdd 17_16/OEN 17_16/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1405 17_16/a_62_902# 17_16/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1406 17_16/a_62_82# 17_16/a_58_538# 17_16/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1407 Vdd 17_16/DATA 17_16/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1408 Vdd 17_16/DIB 17_16/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1409 17_16/DATA 17_16/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1410 GND 17_27/DO 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1411 GND 17_27/a_26_538# 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1412 17_27/DATA 17_27/a_420_786# 17_27/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1413 17_27/DIB 17_27/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1414 17_27/a_62_902# 17_27/a_26_538# 17_27/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1415 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1416 17_27/DI 17_27/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1417 Vdd 17_27/DO 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1418 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1419 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1420 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1421 Vdd 17_27/a_58_538# 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1422 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1423 GND 17_27/a_26_538# 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1424 17_27/a_62_902# 17_27/a_58_538# 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1425 17_27/DIB 17_27/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1426 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1427 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1428 17_27/a_62_82# 17_27/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1429 17_27/DI 17_27/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1430 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1431 17_27/a_62_82# 17_27/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1432 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1433 17_27/DATA 17_27/a_252_786# 17_27/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1434 Vdd 17_27/a_58_538# 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1435 17_27/a_62_82# 17_27/a_26_538# 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1436 GND 17_27/DATA 17_27/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1437 GND 17_27/DIB 17_27/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1438 17_27/a_62_902# 17_27/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1439 17_27/a_62_902# 17_27/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1440 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1441 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1442 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1443 17_27/a_62_82# 17_27/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1444 17_27/a_62_82# 17_27/a_58_538# 17_27/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1445 Vdd 17_27/DATA 17_27/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1446 Vdd 17_27/DIB 17_27/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1447 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1448 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1449 17_27/a_62_902# 17_27/a_26_538# 17_27/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1450 17_27/DIB 17_27/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1451 17_27/DI 17_27/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1452 17_27/a_62_902# 17_27/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1453 GND 17_27/DO 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1454 GND 17_27/DO 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1455 17_27/a_58_538# 17_27/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1456 17_27/a_62_902# 17_27/a_58_538# 17_27/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1457 17_27/DI 17_27/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1458 Vdd 17_27/DO 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1459 17_27/DIB 17_27/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1460 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1461 17_27/DIB 17_27/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1462 17_27/DI 17_27/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1463 GND 17_27/DATA 17_27/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1464 17_27/a_58_538# 17_27/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1465 Vdd 17_27/DO 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1466 17_27/a_62_82# 17_27/a_26_538# 17_27/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1467 GND 17_27/DIB 17_27/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1468 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1469 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1470 17_27/DIB 17_27/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1471 17_27/DI 17_27/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1472 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1473 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1474 17_27/a_62_82# 17_27/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1475 GND 17_27/a_62_82# 17_27/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1476 GND 17_27/OEN 17_27/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1477 17_27/a_62_82# 17_27/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1478 Vdd 17_27/DATA 17_27/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1479 Vdd 17_27/DIB 17_27/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1480 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1481 17_27/DATA 17_27/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1482 Vdd 17_27/a_62_902# 17_27/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1483 GND 17_27/DATA 17_27/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1484 GND 17_27/DIB 17_27/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1485 17_27/a_62_902# 17_27/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1486 Vdd 17_27/OEN 17_27/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1487 17_27/a_62_902# 17_27/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1488 17_27/a_62_82# 17_27/a_58_538# 17_27/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1489 Vdd 17_27/DATA 17_27/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1490 Vdd 17_27/DIB 17_27/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1491 17_27/DATA 17_27/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1492 GND 17_17/DO 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1493 GND 17_17/a_26_538# 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1494 17_17/DATA 17_17/a_420_786# 17_17/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1495 17_17/DIB 17_17/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1496 17_17/a_62_902# 17_17/a_26_538# 17_17/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1497 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1498 17_17/DI 17_17/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1499 Vdd 17_17/DO 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1500 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1501 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1502 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1503 Vdd 17_17/a_58_538# 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1504 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1505 GND 17_17/a_26_538# 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1506 17_17/a_62_902# 17_17/a_58_538# 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1507 17_17/DIB 17_17/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1508 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1509 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1510 17_17/a_62_82# 17_17/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1511 17_17/DI 17_17/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1512 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1513 17_17/a_62_82# 17_17/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1514 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1515 17_17/DATA 17_17/a_252_786# 17_17/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1516 Vdd 17_17/a_58_538# 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1517 17_17/a_62_82# 17_17/a_26_538# 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1518 GND 17_17/DATA 17_17/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1519 GND 17_17/DIB 17_17/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1520 17_17/a_62_902# 17_17/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1521 17_17/a_62_902# 17_17/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1522 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1523 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1524 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1525 17_17/a_62_82# 17_17/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1526 17_17/a_62_82# 17_17/a_58_538# 17_17/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1527 Vdd 17_17/DATA 17_17/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1528 Vdd 17_17/DIB 17_17/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1529 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1530 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1531 17_17/a_62_902# 17_17/a_26_538# 17_17/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1532 17_17/DIB 17_17/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1533 17_17/DI 17_17/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1534 17_17/a_62_902# 17_17/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1535 GND 17_17/DO 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1536 GND 17_17/DO 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1537 17_17/a_58_538# 17_17/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1538 17_17/a_62_902# 17_17/a_58_538# 17_17/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1539 17_17/DI 17_17/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1540 Vdd 17_17/DO 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1541 17_17/DIB 17_17/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1542 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1543 17_17/DIB 17_17/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1544 17_17/DI 17_17/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1545 GND 17_17/DATA 17_17/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1546 17_17/a_58_538# 17_17/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1547 Vdd 17_17/DO 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1548 17_17/a_62_82# 17_17/a_26_538# 17_17/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1549 GND 17_17/DIB 17_17/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1550 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1551 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1552 17_17/DIB 17_17/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1553 17_17/DI 17_17/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1554 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1555 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1556 17_17/a_62_82# 17_17/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1557 GND 17_17/a_62_82# 17_17/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1558 GND 17_17/OEN 17_17/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1559 17_17/a_62_82# 17_17/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1560 Vdd 17_17/DATA 17_17/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1561 Vdd 17_17/DIB 17_17/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1562 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1563 17_17/DATA 17_17/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1564 Vdd 17_17/a_62_902# 17_17/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1565 GND 17_17/DATA 17_17/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1566 GND 17_17/DIB 17_17/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1567 17_17/a_62_902# 17_17/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1568 Vdd 17_17/OEN 17_17/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1569 17_17/a_62_902# 17_17/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1570 17_17/a_62_82# 17_17/a_58_538# 17_17/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1571 Vdd 17_17/DATA 17_17/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1572 Vdd 17_17/DIB 17_17/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1573 17_17/DATA 17_17/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1574 GND 17_28/DO 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1575 GND 17_28/a_26_538# 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1576 17_28/DATA 17_28/a_420_786# 17_28/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1577 17_28/DIB 17_28/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1578 17_28/a_62_902# 17_28/a_26_538# 17_28/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1579 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1580 17_28/DI 17_28/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1581 Vdd 17_28/DO 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1582 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1583 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1584 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1585 Vdd 17_28/a_58_538# 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1586 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1587 GND 17_28/a_26_538# 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1588 17_28/a_62_902# 17_28/a_58_538# 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1589 17_28/DIB 17_28/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1590 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1591 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1592 17_28/a_62_82# 17_28/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1593 17_28/DI 17_28/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1594 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1595 17_28/a_62_82# 17_28/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1596 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1597 17_28/DATA 17_28/a_252_786# 17_28/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1598 Vdd 17_28/a_58_538# 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1599 17_28/a_62_82# 17_28/a_26_538# 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1600 GND 17_28/DATA 17_28/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1601 GND 17_28/DIB 17_28/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1602 17_28/a_62_902# 17_28/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1603 17_28/a_62_902# 17_28/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1604 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1605 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1606 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1607 17_28/a_62_82# 17_28/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1608 17_28/a_62_82# 17_28/a_58_538# 17_28/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1609 Vdd 17_28/DATA 17_28/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1610 Vdd 17_28/DIB 17_28/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1611 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1612 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1613 17_28/a_62_902# 17_28/a_26_538# 17_28/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1614 17_28/DIB 17_28/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1615 17_28/DI 17_28/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1616 17_28/a_62_902# 17_28/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1617 GND 17_28/DO 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1618 GND 17_28/DO 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1619 17_28/a_58_538# 17_28/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1620 17_28/a_62_902# 17_28/a_58_538# 17_28/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1621 17_28/DI 17_28/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1622 Vdd 17_28/DO 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1623 17_28/DIB 17_28/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1624 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1625 17_28/DIB 17_28/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1626 17_28/DI 17_28/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1627 GND 17_28/DATA 17_28/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1628 17_28/a_58_538# 17_28/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1629 Vdd 17_28/DO 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1630 17_28/a_62_82# 17_28/a_26_538# 17_28/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1631 GND 17_28/DIB 17_28/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1632 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1633 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1634 17_28/DIB 17_28/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1635 17_28/DI 17_28/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1636 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1637 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1638 17_28/a_62_82# 17_28/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1639 GND 17_28/a_62_82# 17_28/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1640 GND 17_28/OEN 17_28/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1641 17_28/a_62_82# 17_28/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1642 Vdd 17_28/DATA 17_28/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1643 Vdd 17_28/DIB 17_28/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1644 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1645 17_28/DATA 17_28/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1646 Vdd 17_28/a_62_902# 17_28/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1647 GND 17_28/DATA 17_28/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1648 GND 17_28/DIB 17_28/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1649 17_28/a_62_902# 17_28/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1650 Vdd 17_28/OEN 17_28/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1651 17_28/a_62_902# 17_28/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1652 17_28/a_62_82# 17_28/a_58_538# 17_28/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1653 Vdd 17_28/DATA 17_28/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1654 Vdd 17_28/DIB 17_28/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1655 17_28/DATA 17_28/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1656 GND 17_18/DO 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1657 GND 17_18/a_26_538# 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1658 17_18/DATA 17_18/a_420_786# 17_18/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1659 17_18/DIB 17_18/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1660 17_18/a_62_902# 17_18/a_26_538# 17_18/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1661 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1662 17_18/DI 17_18/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1663 Vdd 17_18/DO 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1664 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1665 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1666 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1667 Vdd 17_18/a_58_538# 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1668 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1669 GND 17_18/a_26_538# 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1670 17_18/a_62_902# 17_18/a_58_538# 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1671 17_18/DIB 17_18/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1672 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1673 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1674 17_18/a_62_82# 17_18/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1675 17_18/DI 17_18/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1676 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1677 17_18/a_62_82# 17_18/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1678 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1679 17_18/DATA 17_18/a_252_786# 17_18/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1680 Vdd 17_18/a_58_538# 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1681 17_18/a_62_82# 17_18/a_26_538# 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1682 GND 17_18/DATA 17_18/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1683 GND 17_18/DIB 17_18/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1684 17_18/a_62_902# 17_18/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1685 17_18/a_62_902# 17_18/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1686 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1687 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1688 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1689 17_18/a_62_82# 17_18/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1690 17_18/a_62_82# 17_18/a_58_538# 17_18/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1691 Vdd 17_18/DATA 17_18/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1692 Vdd 17_18/DIB 17_18/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1693 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1694 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1695 17_18/a_62_902# 17_18/a_26_538# 17_18/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1696 17_18/DIB 17_18/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1697 17_18/DI 17_18/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1698 17_18/a_62_902# 17_18/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1699 GND 17_18/DO 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1700 GND 17_18/DO 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1701 17_18/a_58_538# 17_18/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1702 17_18/a_62_902# 17_18/a_58_538# 17_18/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1703 17_18/DI 17_18/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1704 Vdd 17_18/DO 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1705 17_18/DIB 17_18/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1706 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1707 17_18/DIB 17_18/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1708 17_18/DI 17_18/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1709 GND 17_18/DATA 17_18/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1710 17_18/a_58_538# 17_18/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1711 Vdd 17_18/DO 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1712 17_18/a_62_82# 17_18/a_26_538# 17_18/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1713 GND 17_18/DIB 17_18/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1714 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1715 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1716 17_18/DIB 17_18/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1717 17_18/DI 17_18/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1718 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1719 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1720 17_18/a_62_82# 17_18/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1721 GND 17_18/a_62_82# 17_18/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1722 GND 17_18/OEN 17_18/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1723 17_18/a_62_82# 17_18/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1724 Vdd 17_18/DATA 17_18/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1725 Vdd 17_18/DIB 17_18/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1726 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1727 17_18/DATA 17_18/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1728 Vdd 17_18/a_62_902# 17_18/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1729 GND 17_18/DATA 17_18/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1730 GND 17_18/DIB 17_18/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1731 17_18/a_62_902# 17_18/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1732 Vdd 17_18/OEN 17_18/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1733 17_18/a_62_902# 17_18/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1734 17_18/a_62_82# 17_18/a_58_538# 17_18/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1735 Vdd 17_18/DATA 17_18/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1736 Vdd 17_18/DIB 17_18/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1737 17_18/DATA 17_18/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1738 i b GND Gnd nfet w=20 l=4
+  ad=0.12n pd=32u as=0.2n ps=60u
M1739 i a hwtest_0/NOR2X1_0/a_18_108# Vdd pfet w=80 l=4
+  ad=0.8n pd=0.18m as=0.24n ps=86u
M1740 GND a i Gnd nfet w=20 l=4
+  ad=0.2n pd=60u as=0.12n ps=32u
M1741 hwtest_0/NOR2X1_0/a_18_108# b Vdd Vdd pfet w=80 l=4
+  ad=0.24n pd=86u as=0.8n ps=0.18m
M1742 hwtest_0/NOR2X1_1/Y d GND Gnd nfet w=20 l=4
+  ad=0.24n pd=64u as=0 ps=0
M1743 hwtest_0/NOR2X1_1/Y i hwtest_0/NOR2X1_1/a_18_108# Vdd pfet w=80 l=4
+  ad=0.8n pd=0.18m as=0.48n ps=0.172m
M1744 GND i hwtest_0/NOR2X1_1/Y Gnd nfet w=20 l=4
+  ad=0 pd=0 as=0 ps=0
M1745 hwtest_0/NOR2X1_1/a_18_108# d Vdd Vdd pfet w=80 l=4
+  ad=0 pd=0 as=0 ps=0
M1746 h hwtest_0/AND2X2_0/a_4_12# GND Gnd nfet w=40 l=4
+  ad=0.4n pd=100u as=0.24n ps=52u
M1747 hwtest_0/AND2X2_0/a_18_12# hwtest_0/NOR2X1_1/Y hwtest_0/AND2X2_0/a_4_12# Gnd nfet w=40 l=4
+  ad=0.12n pd=46u as=0.4n ps=100u
M1748 Vdd c hwtest_0/AND2X2_0/a_4_12# Vdd pfet w=40 l=4
+  ad=0.432n pd=92u as=0.24n ps=52u
M1749 h hwtest_0/AND2X2_0/a_4_12# Vdd Vdd pfet w=80 l=4
+  ad=0.8n pd=0.18m as=0.432n ps=92u
M1750 GND c hwtest_0/AND2X2_0/a_18_12# Gnd nfet w=40 l=4
+  ad=0.24n pd=52u as=0.12n ps=46u
M1751 hwtest_0/AND2X2_0/a_4_12# hwtest_0/NOR2X1_1/Y Vdd Vdd pfet w=40 l=4
+  ad=0.24n pd=52u as=0.4n ps=100u
M1752 GND 17_29/DO 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1753 GND 17_29/a_26_538# 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1754 17_29/DATA 17_29/a_420_786# 17_29/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1755 17_29/DIB 17_29/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1756 17_29/a_62_902# 17_29/a_26_538# 17_29/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1757 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1758 17_29/DI 17_29/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1759 Vdd 17_29/DO 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1760 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1761 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1762 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1763 Vdd 17_29/a_58_538# 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1764 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1765 GND 17_29/a_26_538# 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1766 17_29/a_62_902# 17_29/a_58_538# 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1767 17_29/DIB 17_29/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1768 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1769 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1770 17_29/a_62_82# 17_29/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1771 17_29/DI 17_29/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1772 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1773 17_29/a_62_82# 17_29/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1774 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1775 17_29/DATA 17_29/a_252_786# 17_29/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1776 Vdd 17_29/a_58_538# 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1777 17_29/a_62_82# 17_29/a_26_538# 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1778 GND 17_29/DATA 17_29/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1779 GND 17_29/DIB 17_29/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1780 17_29/a_62_902# 17_29/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1781 17_29/a_62_902# 17_29/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1782 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1783 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1784 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1785 17_29/a_62_82# 17_29/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1786 17_29/a_62_82# 17_29/a_58_538# 17_29/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1787 Vdd 17_29/DATA 17_29/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1788 Vdd 17_29/DIB 17_29/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1789 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1790 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1791 17_29/a_62_902# 17_29/a_26_538# 17_29/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1792 17_29/DIB 17_29/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1793 17_29/DI 17_29/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1794 17_29/a_62_902# 17_29/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1795 GND 17_29/DO 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1796 GND 17_29/DO 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1797 17_29/a_58_538# 17_29/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1798 17_29/a_62_902# 17_29/a_58_538# 17_29/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1799 17_29/DI 17_29/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1800 Vdd 17_29/DO 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1801 17_29/DIB 17_29/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1802 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1803 17_29/DIB 17_29/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1804 17_29/DI 17_29/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1805 GND 17_29/DATA 17_29/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1806 17_29/a_58_538# 17_29/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1807 Vdd 17_29/DO 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1808 17_29/a_62_82# 17_29/a_26_538# 17_29/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1809 GND 17_29/DIB 17_29/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1810 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1811 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1812 17_29/DIB 17_29/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1813 17_29/DI 17_29/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1814 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1815 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1816 17_29/a_62_82# 17_29/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1817 GND 17_29/a_62_82# 17_29/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1818 GND 17_29/OEN 17_29/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1819 17_29/a_62_82# 17_29/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1820 Vdd 17_29/DATA 17_29/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1821 Vdd 17_29/DIB 17_29/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1822 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1823 17_29/DATA 17_29/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1824 Vdd 17_29/a_62_902# 17_29/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1825 GND 17_29/DATA 17_29/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1826 GND 17_29/DIB 17_29/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1827 17_29/a_62_902# 17_29/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1828 Vdd 17_29/OEN 17_29/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1829 17_29/a_62_902# 17_29/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1830 17_29/a_62_82# 17_29/a_58_538# 17_29/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1831 Vdd 17_29/DATA 17_29/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1832 Vdd 17_29/DIB 17_29/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1833 17_29/DATA 17_29/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1834 GND 17_19/DO 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1835 GND 17_19/a_26_538# 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1836 17_19/DATA 17_19/a_420_786# 17_19/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1837 17_19/DIB 17_19/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1838 17_19/a_62_902# 17_19/a_26_538# 17_19/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1839 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1840 17_19/DI 17_19/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1841 Vdd 17_19/DO 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1842 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1843 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1844 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1845 Vdd 17_19/a_58_538# 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1846 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1847 GND 17_19/a_26_538# 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1848 17_19/a_62_902# 17_19/a_58_538# 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1849 17_19/DIB 17_19/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1850 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1851 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1852 17_19/a_62_82# 17_19/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1853 17_19/DI 17_19/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1854 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1855 17_19/a_62_82# 17_19/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1856 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1857 17_19/DATA 17_19/a_252_786# 17_19/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1858 Vdd 17_19/a_58_538# 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1859 17_19/a_62_82# 17_19/a_26_538# 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1860 GND 17_19/DATA 17_19/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1861 GND 17_19/DIB 17_19/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1862 17_19/a_62_902# 17_19/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1863 17_19/a_62_902# 17_19/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1864 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1865 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1866 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1867 17_19/a_62_82# 17_19/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1868 17_19/a_62_82# 17_19/a_58_538# 17_19/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1869 Vdd 17_19/DATA 17_19/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1870 Vdd 17_19/DIB 17_19/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1871 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1872 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1873 17_19/a_62_902# 17_19/a_26_538# 17_19/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1874 17_19/DIB 17_19/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1875 17_19/DI 17_19/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1876 17_19/a_62_902# 17_19/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1877 GND 17_19/DO 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1878 GND 17_19/DO 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1879 17_19/a_58_538# 17_19/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1880 17_19/a_62_902# 17_19/a_58_538# 17_19/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1881 17_19/DI 17_19/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1882 Vdd 17_19/DO 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1883 17_19/DIB 17_19/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1884 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1885 17_19/DIB 17_19/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1886 17_19/DI 17_19/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1887 GND 17_19/DATA 17_19/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1888 17_19/a_58_538# 17_19/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1889 Vdd 17_19/DO 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1890 17_19/a_62_82# 17_19/a_26_538# 17_19/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1891 GND 17_19/DIB 17_19/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1892 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1893 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1894 17_19/DIB 17_19/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1895 17_19/DI 17_19/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1896 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1897 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1898 17_19/a_62_82# 17_19/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1899 GND 17_19/a_62_82# 17_19/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1900 GND 17_19/OEN 17_19/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M1901 17_19/a_62_82# 17_19/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1902 Vdd 17_19/DATA 17_19/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1903 Vdd 17_19/DIB 17_19/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1904 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1905 17_19/DATA 17_19/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1906 Vdd 17_19/a_62_902# 17_19/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1907 GND 17_19/DATA 17_19/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1908 GND 17_19/DIB 17_19/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1909 17_19/a_62_902# 17_19/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1910 Vdd 17_19/OEN 17_19/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M1911 17_19/a_62_902# 17_19/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1912 17_19/a_62_82# 17_19/a_58_538# 17_19/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1913 Vdd 17_19/DATA 17_19/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1914 Vdd 17_19/DIB 17_19/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1915 17_19/DATA 17_19/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1916 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1917 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1918 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.4n ps=0.234m
M1919 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M1920 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.4n pd=0.234m as=8.2n ps=0.282m
M1921 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M1922 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.2n ps=0.282m
M1923 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M1924 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.4n ps=0.234m
M1925 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M1926 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.4n pd=0.234m as=8.2n ps=0.282m
M1927 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.2n ps=0.282m
M1928 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=11.328096u ps=0.41559
M1929 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1930 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1931 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1932 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1933 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1934 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1935 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1936 GND Vdd Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1937 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1938 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1939 Vdd Vdd GND Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1940 GND 17_1/DO 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M1941 GND 17_1/a_26_538# 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1942 17_1/DATA 17_1/a_420_786# 17_1/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M1943 17_1/DIB 17_1/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1944 17_1/a_62_902# 17_1/a_26_538# 17_1/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M1945 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M1946 17_1/DI 17_1/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M1947 Vdd 17_1/DO 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1948 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M1949 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1950 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1951 Vdd 17_1/a_58_538# 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1952 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1953 GND 17_1/a_26_538# 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1954 17_1/a_62_902# 17_1/a_58_538# 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M1955 17_1/DIB 17_1/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1956 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1957 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1958 17_1/a_62_82# 17_1/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1959 17_1/DI 17_1/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M1960 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1961 17_1/a_62_82# 17_1/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1962 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1963 17_1/DATA 17_1/a_252_786# 17_1/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M1964 Vdd 17_1/a_58_538# 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1965 17_1/a_62_82# 17_1/a_26_538# 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1966 GND 17_1/DATA 17_1/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1967 GND 17_1/DIB 17_1/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1968 17_1/a_62_902# 17_1/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1969 17_1/a_62_902# 17_1/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1970 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1971 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1972 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1973 17_1/a_62_82# 17_1/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1974 17_1/a_62_82# 17_1/a_58_538# 17_1/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1975 Vdd 17_1/DATA 17_1/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1976 Vdd 17_1/DIB 17_1/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1977 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1978 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1979 17_1/a_62_902# 17_1/a_26_538# 17_1/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1980 17_1/DIB 17_1/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1981 17_1/DI 17_1/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1982 17_1/a_62_902# 17_1/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1983 GND 17_1/DO 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1984 GND 17_1/DO 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1985 17_1/a_58_538# 17_1/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M1986 17_1/a_62_902# 17_1/a_58_538# 17_1/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1987 17_1/DI 17_1/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1988 Vdd 17_1/DO 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1989 17_1/DIB 17_1/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1990 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1991 17_1/DIB 17_1/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1992 17_1/DI 17_1/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1993 GND 17_1/DATA 17_1/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1994 17_1/a_58_538# 17_1/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M1995 Vdd 17_1/DO 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1996 17_1/a_62_82# 17_1/a_26_538# 17_1/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M1997 GND 17_1/DIB 17_1/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M1998 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M1999 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2000 17_1/DIB 17_1/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2001 17_1/DI 17_1/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2002 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2003 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2004 17_1/a_62_82# 17_1/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2005 GND 17_1/a_62_82# 17_1/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2006 GND 17_1/OEN 17_1/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2007 17_1/a_62_82# 17_1/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2008 Vdd 17_1/DATA 17_1/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2009 Vdd 17_1/DIB 17_1/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2010 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2011 17_1/DATA 17_1/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2012 Vdd 17_1/a_62_902# 17_1/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2013 GND 17_1/DATA 17_1/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2014 GND 17_1/DIB 17_1/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2015 17_1/a_62_902# 17_1/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2016 Vdd 17_1/OEN 17_1/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2017 17_1/a_62_902# 17_1/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2018 17_1/a_62_82# 17_1/a_58_538# 17_1/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2019 Vdd 17_1/DATA 17_1/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2020 Vdd 17_1/DIB 17_1/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2021 17_1/DATA 17_1/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2022 GND 17_0/DO 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2023 GND 17_0/a_26_538# 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2024 17_0/DATA 17_0/a_420_786# 17_0/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2025 17_0/DIB 17_0/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2026 17_0/a_62_902# 17_0/a_26_538# 17_0/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2027 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2028 17_0/DI 17_0/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2029 Vdd 17_0/DO 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2030 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2031 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2032 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2033 Vdd 17_0/a_58_538# 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2034 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2035 GND 17_0/a_26_538# 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2036 17_0/a_62_902# 17_0/a_58_538# 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2037 17_0/DIB 17_0/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2038 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2039 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2040 17_0/a_62_82# 17_0/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2041 17_0/DI 17_0/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2042 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2043 17_0/a_62_82# 17_0/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2044 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2045 17_0/DATA 17_0/a_252_786# 17_0/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2046 Vdd 17_0/a_58_538# 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2047 17_0/a_62_82# 17_0/a_26_538# 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2048 GND 17_0/DATA 17_0/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2049 GND 17_0/DIB 17_0/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2050 17_0/a_62_902# 17_0/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2051 17_0/a_62_902# 17_0/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2052 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2053 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2054 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2055 17_0/a_62_82# 17_0/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2056 17_0/a_62_82# 17_0/a_58_538# 17_0/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2057 Vdd 17_0/DATA 17_0/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2058 Vdd 17_0/DIB 17_0/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2059 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2060 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2061 17_0/a_62_902# 17_0/a_26_538# 17_0/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2062 17_0/DIB 17_0/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2063 17_0/DI 17_0/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2064 17_0/a_62_902# 17_0/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2065 GND 17_0/DO 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2066 GND 17_0/DO 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2067 17_0/a_58_538# 17_0/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2068 17_0/a_62_902# 17_0/a_58_538# 17_0/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2069 17_0/DI 17_0/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2070 Vdd 17_0/DO 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2071 17_0/DIB 17_0/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2072 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2073 17_0/DIB 17_0/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2074 17_0/DI 17_0/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2075 GND 17_0/DATA 17_0/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2076 17_0/a_58_538# 17_0/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2077 Vdd 17_0/DO 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2078 17_0/a_62_82# 17_0/a_26_538# 17_0/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2079 GND 17_0/DIB 17_0/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2080 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2081 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2082 17_0/DIB 17_0/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2083 17_0/DI 17_0/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2084 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2085 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2086 17_0/a_62_82# 17_0/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2087 GND 17_0/a_62_82# 17_0/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2088 GND GND 17_0/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2089 17_0/a_62_82# 17_0/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2090 Vdd 17_0/DATA 17_0/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2091 Vdd 17_0/DIB 17_0/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2092 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2093 17_0/DATA 17_0/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2094 Vdd 17_0/a_62_902# 17_0/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2095 GND 17_0/DATA 17_0/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2096 GND 17_0/DIB 17_0/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2097 17_0/a_62_902# 17_0/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2098 Vdd GND 17_0/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2099 17_0/a_62_902# 17_0/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2100 17_0/a_62_82# 17_0/a_58_538# 17_0/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2101 Vdd 17_0/DATA 17_0/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2102 Vdd 17_0/DIB 17_0/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2103 17_0/DATA 17_0/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2104 GND 17_2/DO 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2105 GND 17_2/a_26_538# 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2106 p_a 17_2/a_420_786# p_a Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2107 17_2/DIB p_a GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2108 17_2/a_62_902# 17_2/a_26_538# 17_2/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2109 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2110 a 17_2/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2111 Vdd 17_2/DO 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2112 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2113 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2114 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2115 Vdd 17_2/a_58_538# 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2116 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2117 GND 17_2/a_26_538# 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2118 17_2/a_62_902# 17_2/a_58_538# 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2119 17_2/DIB p_a Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2120 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2121 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2122 17_2/a_62_82# 17_2/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2123 a 17_2/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2124 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2125 17_2/a_62_82# 17_2/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2126 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2127 p_a 17_2/a_252_786# p_a Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2128 Vdd 17_2/a_58_538# 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2129 17_2/a_62_82# 17_2/a_26_538# 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2130 GND p_a 17_2/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2131 GND 17_2/DIB a Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2132 17_2/a_62_902# 17_2/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2133 17_2/a_62_902# 17_2/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2134 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2135 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2136 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2137 17_2/a_62_82# 17_2/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2138 17_2/a_62_82# 17_2/a_58_538# 17_2/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2139 Vdd p_a 17_2/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2140 Vdd 17_2/DIB a Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2141 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2142 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2143 17_2/a_62_902# 17_2/a_26_538# 17_2/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2144 17_2/DIB p_a GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2145 a 17_2/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2146 17_2/a_62_902# 17_2/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2147 GND 17_2/DO 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2148 GND 17_2/DO 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2149 17_2/a_58_538# 17_2/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2150 17_2/a_62_902# 17_2/a_58_538# 17_2/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2151 a 17_2/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2152 Vdd 17_2/DO 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2153 17_2/DIB p_a Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2154 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2155 17_2/DIB p_a GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2156 a 17_2/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2157 GND p_a 17_2/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2158 17_2/a_58_538# 17_2/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2159 Vdd 17_2/DO 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2160 17_2/a_62_82# 17_2/a_26_538# 17_2/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2161 GND 17_2/DIB a Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2162 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2163 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2164 17_2/DIB p_a Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2165 a 17_2/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2166 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2167 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2168 17_2/a_62_82# 17_2/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2169 GND 17_2/a_62_82# p_a GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2170 GND GND 17_2/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2171 17_2/a_62_82# 17_2/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2172 Vdd p_a 17_2/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2173 Vdd 17_2/DIB a Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2174 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2175 p_a 17_2/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2176 Vdd 17_2/a_62_902# p_a Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2177 GND p_a 17_2/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2178 GND 17_2/DIB a Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2179 17_2/a_62_902# 17_2/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2180 Vdd GND 17_2/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2181 17_2/a_62_902# 17_2/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2182 17_2/a_62_82# 17_2/a_58_538# 17_2/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2183 Vdd p_a 17_2/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2184 Vdd 17_2/DIB a Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2185 p_a 17_2/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2186 GND i 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2187 GND 17_3/a_26_538# 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2188 p_i 17_3/a_420_786# p_i Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2189 17_3/DIB p_i GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2190 17_3/a_62_902# 17_3/a_26_538# 17_3/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2191 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2192 17_3/DI 17_3/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2193 Vdd i 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2194 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2195 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2196 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2197 Vdd 17_3/a_58_538# 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2198 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2199 GND 17_3/a_26_538# 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2200 17_3/a_62_902# 17_3/a_58_538# 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2201 17_3/DIB p_i Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2202 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2203 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2204 17_3/a_62_82# 17_3/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2205 17_3/DI 17_3/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2206 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2207 17_3/a_62_82# i GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2208 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2209 p_i 17_3/a_252_786# p_i Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2210 Vdd 17_3/a_58_538# 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2211 17_3/a_62_82# 17_3/a_26_538# 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2212 GND p_i 17_3/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2213 GND 17_3/DIB 17_3/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2214 17_3/a_62_902# 17_3/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2215 17_3/a_62_902# i Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2216 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2217 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2218 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2219 17_3/a_62_82# 17_3/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2220 17_3/a_62_82# 17_3/a_58_538# 17_3/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2221 Vdd p_i 17_3/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2222 Vdd 17_3/DIB 17_3/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2223 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2224 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2225 17_3/a_62_902# 17_3/a_26_538# 17_3/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2226 17_3/DIB p_i GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2227 17_3/DI 17_3/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2228 17_3/a_62_902# 17_3/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2229 GND i 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2230 GND i 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2231 17_3/a_58_538# 17_3/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2232 17_3/a_62_902# 17_3/a_58_538# 17_3/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2233 17_3/DI 17_3/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2234 Vdd i 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2235 17_3/DIB p_i Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2236 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2237 17_3/DIB p_i GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2238 17_3/DI 17_3/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2239 GND p_i 17_3/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2240 17_3/a_58_538# 17_3/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2241 Vdd i 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2242 17_3/a_62_82# 17_3/a_26_538# 17_3/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2243 GND 17_3/DIB 17_3/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2244 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2245 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2246 17_3/DIB p_i Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2247 17_3/DI 17_3/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2248 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2249 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2250 17_3/a_62_82# 17_3/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2251 GND 17_3/a_62_82# p_i GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2252 GND Vdd 17_3/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2253 17_3/a_62_82# i GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2254 Vdd p_i 17_3/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2255 Vdd 17_3/DIB 17_3/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2256 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2257 p_i 17_3/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2258 Vdd 17_3/a_62_902# p_i Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2259 GND p_i 17_3/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2260 GND 17_3/DIB 17_3/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2261 17_3/a_62_902# 17_3/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2262 Vdd Vdd 17_3/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2263 17_3/a_62_902# i Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2264 17_3/a_62_82# 17_3/a_58_538# 17_3/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2265 Vdd p_i 17_3/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2266 Vdd 17_3/DIB 17_3/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2267 p_i 17_3/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2268 GND 17_4/DO 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2269 GND 17_4/a_26_538# 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2270 p_b 17_4/a_420_786# p_b Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2271 17_4/DIB p_b GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2272 17_4/a_62_902# 17_4/a_26_538# 17_4/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2273 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2274 b 17_4/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2275 Vdd 17_4/DO 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2276 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2277 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2278 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2279 Vdd 17_4/a_58_538# 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2280 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2281 GND 17_4/a_26_538# 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2282 17_4/a_62_902# 17_4/a_58_538# 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2283 17_4/DIB p_b Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2284 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2285 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2286 17_4/a_62_82# 17_4/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2287 b 17_4/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2288 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2289 17_4/a_62_82# 17_4/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2290 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2291 p_b 17_4/a_252_786# p_b Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2292 Vdd 17_4/a_58_538# 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2293 17_4/a_62_82# 17_4/a_26_538# 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2294 GND p_b 17_4/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2295 GND 17_4/DIB b Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2296 17_4/a_62_902# 17_4/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2297 17_4/a_62_902# 17_4/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2298 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2299 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2300 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2301 17_4/a_62_82# 17_4/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2302 17_4/a_62_82# 17_4/a_58_538# 17_4/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2303 Vdd p_b 17_4/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2304 Vdd 17_4/DIB b Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2305 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2306 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2307 17_4/a_62_902# 17_4/a_26_538# 17_4/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2308 17_4/DIB p_b GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2309 b 17_4/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2310 17_4/a_62_902# 17_4/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2311 GND 17_4/DO 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2312 GND 17_4/DO 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2313 17_4/a_58_538# 17_4/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2314 17_4/a_62_902# 17_4/a_58_538# 17_4/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2315 b 17_4/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2316 Vdd 17_4/DO 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2317 17_4/DIB p_b Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2318 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2319 17_4/DIB p_b GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2320 b 17_4/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2321 GND p_b 17_4/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2322 17_4/a_58_538# 17_4/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2323 Vdd 17_4/DO 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2324 17_4/a_62_82# 17_4/a_26_538# 17_4/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2325 GND 17_4/DIB b Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2326 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2327 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2328 17_4/DIB p_b Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2329 b 17_4/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2330 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2331 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2332 17_4/a_62_82# 17_4/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2333 GND 17_4/a_62_82# p_b GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2334 GND GND 17_4/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2335 17_4/a_62_82# 17_4/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2336 Vdd p_b 17_4/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2337 Vdd 17_4/DIB b Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2338 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2339 p_b 17_4/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2340 Vdd 17_4/a_62_902# p_b Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2341 GND p_b 17_4/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2342 GND 17_4/DIB b Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2343 17_4/a_62_902# 17_4/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2344 Vdd GND 17_4/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2345 17_4/a_62_902# 17_4/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2346 17_4/a_62_82# 17_4/a_58_538# 17_4/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2347 Vdd p_b 17_4/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2348 Vdd 17_4/DIB b Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2349 p_b 17_4/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2350 GND 17_5/DO 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2351 GND 17_5/a_26_538# 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2352 p_d 17_5/a_420_786# p_d Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2353 17_5/DIB p_d GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2354 17_5/a_62_902# 17_5/a_26_538# 17_5/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2355 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2356 d 17_5/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2357 Vdd 17_5/DO 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2358 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2359 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2360 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2361 Vdd 17_5/a_58_538# 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2362 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2363 GND 17_5/a_26_538# 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2364 17_5/a_62_902# 17_5/a_58_538# 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2365 17_5/DIB p_d Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2366 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2367 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2368 17_5/a_62_82# 17_5/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2369 d 17_5/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2370 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2371 17_5/a_62_82# 17_5/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2372 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2373 p_d 17_5/a_252_786# p_d Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2374 Vdd 17_5/a_58_538# 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2375 17_5/a_62_82# 17_5/a_26_538# 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2376 GND p_d 17_5/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2377 GND 17_5/DIB d Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2378 17_5/a_62_902# 17_5/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2379 17_5/a_62_902# 17_5/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2380 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2381 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2382 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2383 17_5/a_62_82# 17_5/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2384 17_5/a_62_82# 17_5/a_58_538# 17_5/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2385 Vdd p_d 17_5/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2386 Vdd 17_5/DIB d Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2387 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2388 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2389 17_5/a_62_902# 17_5/a_26_538# 17_5/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2390 17_5/DIB p_d GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2391 d 17_5/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2392 17_5/a_62_902# 17_5/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2393 GND 17_5/DO 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2394 GND 17_5/DO 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2395 17_5/a_58_538# 17_5/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2396 17_5/a_62_902# 17_5/a_58_538# 17_5/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2397 d 17_5/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2398 Vdd 17_5/DO 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2399 17_5/DIB p_d Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2400 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2401 17_5/DIB p_d GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2402 d 17_5/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2403 GND p_d 17_5/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2404 17_5/a_58_538# 17_5/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2405 Vdd 17_5/DO 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2406 17_5/a_62_82# 17_5/a_26_538# 17_5/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2407 GND 17_5/DIB d Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2408 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2409 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2410 17_5/DIB p_d Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2411 d 17_5/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2412 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2413 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2414 17_5/a_62_82# 17_5/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2415 GND 17_5/a_62_82# p_d GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2416 GND GND 17_5/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2417 17_5/a_62_82# 17_5/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2418 Vdd p_d 17_5/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2419 Vdd 17_5/DIB d Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2420 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2421 p_d 17_5/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2422 Vdd 17_5/a_62_902# p_d Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2423 GND p_d 17_5/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2424 GND 17_5/DIB d Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2425 17_5/a_62_902# 17_5/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2426 Vdd GND 17_5/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2427 17_5/a_62_902# 17_5/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2428 17_5/a_62_82# 17_5/a_58_538# 17_5/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2429 Vdd p_d 17_5/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2430 Vdd 17_5/DIB d Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2431 p_d 17_5/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2432 GND 17_6/DO 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2433 GND 17_6/a_26_538# 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2434 p_c 17_6/a_420_786# p_c Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2435 17_6/DIB p_c GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2436 17_6/a_62_902# 17_6/a_26_538# 17_6/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2437 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2438 c 17_6/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2439 Vdd 17_6/DO 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2440 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2441 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2442 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2443 Vdd 17_6/a_58_538# 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2444 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2445 GND 17_6/a_26_538# 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2446 17_6/a_62_902# 17_6/a_58_538# 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2447 17_6/DIB p_c Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2448 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2449 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2450 17_6/a_62_82# 17_6/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2451 c 17_6/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2452 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2453 17_6/a_62_82# 17_6/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2454 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2455 p_c 17_6/a_252_786# p_c Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2456 Vdd 17_6/a_58_538# 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2457 17_6/a_62_82# 17_6/a_26_538# 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2458 GND p_c 17_6/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2459 GND 17_6/DIB c Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2460 17_6/a_62_902# 17_6/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2461 17_6/a_62_902# 17_6/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2462 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2463 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2464 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2465 17_6/a_62_82# 17_6/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2466 17_6/a_62_82# 17_6/a_58_538# 17_6/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2467 Vdd p_c 17_6/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2468 Vdd 17_6/DIB c Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2469 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2470 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2471 17_6/a_62_902# 17_6/a_26_538# 17_6/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2472 17_6/DIB p_c GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2473 c 17_6/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2474 17_6/a_62_902# 17_6/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2475 GND 17_6/DO 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2476 GND 17_6/DO 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2477 17_6/a_58_538# 17_6/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2478 17_6/a_62_902# 17_6/a_58_538# 17_6/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2479 c 17_6/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2480 Vdd 17_6/DO 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2481 17_6/DIB p_c Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2482 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2483 17_6/DIB p_c GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2484 c 17_6/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2485 GND p_c 17_6/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2486 17_6/a_58_538# 17_6/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2487 Vdd 17_6/DO 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2488 17_6/a_62_82# 17_6/a_26_538# 17_6/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2489 GND 17_6/DIB c Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2490 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2491 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2492 17_6/DIB p_c Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2493 c 17_6/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2494 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2495 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2496 17_6/a_62_82# 17_6/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2497 GND 17_6/a_62_82# p_c GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2498 GND GND 17_6/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2499 17_6/a_62_82# 17_6/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2500 Vdd p_c 17_6/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2501 Vdd 17_6/DIB c Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2502 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2503 p_c 17_6/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2504 Vdd 17_6/a_62_902# p_c Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2505 GND p_c 17_6/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2506 GND 17_6/DIB c Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2507 17_6/a_62_902# 17_6/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2508 Vdd GND 17_6/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2509 17_6/a_62_902# 17_6/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2510 17_6/a_62_82# 17_6/a_58_538# 17_6/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2511 Vdd p_c 17_6/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2512 Vdd 17_6/DIB c Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2513 p_c 17_6/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2514 GND h 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2515 GND 17_7/a_26_538# 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2516 p_h 17_7/a_420_786# p_h Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2517 17_7/DIB p_h GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2518 17_7/a_62_902# 17_7/a_26_538# 17_7/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2519 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2520 17_7/DI 17_7/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2521 Vdd h 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2522 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2523 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2524 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2525 Vdd 17_7/a_58_538# 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2526 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2527 GND 17_7/a_26_538# 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2528 17_7/a_62_902# 17_7/a_58_538# 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2529 17_7/DIB p_h Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2530 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2531 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2532 17_7/a_62_82# 17_7/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2533 17_7/DI 17_7/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2534 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2535 17_7/a_62_82# h GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2536 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2537 p_h 17_7/a_252_786# p_h Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2538 Vdd 17_7/a_58_538# 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2539 17_7/a_62_82# 17_7/a_26_538# 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2540 GND p_h 17_7/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2541 GND 17_7/DIB 17_7/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2542 17_7/a_62_902# 17_7/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2543 17_7/a_62_902# h Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2544 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2545 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2546 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2547 17_7/a_62_82# 17_7/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2548 17_7/a_62_82# 17_7/a_58_538# 17_7/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2549 Vdd p_h 17_7/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2550 Vdd 17_7/DIB 17_7/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2551 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2552 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2553 17_7/a_62_902# 17_7/a_26_538# 17_7/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2554 17_7/DIB p_h GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2555 17_7/DI 17_7/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2556 17_7/a_62_902# 17_7/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2557 GND h 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2558 GND h 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2559 17_7/a_58_538# 17_7/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2560 17_7/a_62_902# 17_7/a_58_538# 17_7/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2561 17_7/DI 17_7/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2562 Vdd h 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2563 17_7/DIB p_h Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2564 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2565 17_7/DIB p_h GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2566 17_7/DI 17_7/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2567 GND p_h 17_7/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2568 17_7/a_58_538# 17_7/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2569 Vdd h 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2570 17_7/a_62_82# 17_7/a_26_538# 17_7/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2571 GND 17_7/DIB 17_7/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2572 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2573 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2574 17_7/DIB p_h Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2575 17_7/DI 17_7/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2576 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2577 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2578 17_7/a_62_82# 17_7/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2579 GND 17_7/a_62_82# p_h GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2580 GND Vdd 17_7/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2581 17_7/a_62_82# h GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2582 Vdd p_h 17_7/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2583 Vdd 17_7/DIB 17_7/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2584 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2585 p_h 17_7/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2586 Vdd 17_7/a_62_902# p_h Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2587 GND p_h 17_7/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2588 GND 17_7/DIB 17_7/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2589 17_7/a_62_902# 17_7/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2590 Vdd Vdd 17_7/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2591 17_7/a_62_902# h Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2592 17_7/a_62_82# 17_7/a_58_538# 17_7/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2593 Vdd p_h 17_7/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2594 Vdd 17_7/DIB 17_7/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2595 p_h 17_7/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2596 GND 17_8/DO 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2597 GND 17_8/a_26_538# 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2598 17_8/DATA 17_8/a_420_786# 17_8/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2599 17_8/DIB 17_8/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2600 17_8/a_62_902# 17_8/a_26_538# 17_8/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2601 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2602 17_8/DI 17_8/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2603 Vdd 17_8/DO 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2604 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2605 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2606 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2607 Vdd 17_8/a_58_538# 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2608 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2609 GND 17_8/a_26_538# 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2610 17_8/a_62_902# 17_8/a_58_538# 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2611 17_8/DIB 17_8/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2612 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2613 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2614 17_8/a_62_82# 17_8/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2615 17_8/DI 17_8/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2616 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2617 17_8/a_62_82# 17_8/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2618 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2619 17_8/DATA 17_8/a_252_786# 17_8/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2620 Vdd 17_8/a_58_538# 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2621 17_8/a_62_82# 17_8/a_26_538# 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2622 GND 17_8/DATA 17_8/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2623 GND 17_8/DIB 17_8/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2624 17_8/a_62_902# 17_8/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2625 17_8/a_62_902# 17_8/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2626 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2627 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2628 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2629 17_8/a_62_82# 17_8/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2630 17_8/a_62_82# 17_8/a_58_538# 17_8/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2631 Vdd 17_8/DATA 17_8/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2632 Vdd 17_8/DIB 17_8/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2633 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2634 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2635 17_8/a_62_902# 17_8/a_26_538# 17_8/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2636 17_8/DIB 17_8/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2637 17_8/DI 17_8/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2638 17_8/a_62_902# 17_8/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2639 GND 17_8/DO 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2640 GND 17_8/DO 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2641 17_8/a_58_538# 17_8/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2642 17_8/a_62_902# 17_8/a_58_538# 17_8/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2643 17_8/DI 17_8/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2644 Vdd 17_8/DO 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2645 17_8/DIB 17_8/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2646 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2647 17_8/DIB 17_8/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2648 17_8/DI 17_8/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2649 GND 17_8/DATA 17_8/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2650 17_8/a_58_538# 17_8/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2651 Vdd 17_8/DO 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2652 17_8/a_62_82# 17_8/a_26_538# 17_8/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2653 GND 17_8/DIB 17_8/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2654 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2655 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2656 17_8/DIB 17_8/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2657 17_8/DI 17_8/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2658 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2659 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2660 17_8/a_62_82# 17_8/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2661 GND 17_8/a_62_82# 17_8/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2662 GND 17_8/OEN 17_8/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2663 17_8/a_62_82# 17_8/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2664 Vdd 17_8/DATA 17_8/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2665 Vdd 17_8/DIB 17_8/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2666 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2667 17_8/DATA 17_8/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2668 Vdd 17_8/a_62_902# 17_8/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2669 GND 17_8/DATA 17_8/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2670 GND 17_8/DIB 17_8/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2671 17_8/a_62_902# 17_8/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2672 Vdd 17_8/OEN 17_8/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2673 17_8/a_62_902# 17_8/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2674 17_8/a_62_82# 17_8/a_58_538# 17_8/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2675 Vdd 17_8/DATA 17_8/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2676 Vdd 17_8/DIB 17_8/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2677 17_8/DATA 17_8/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2678 GND 17_9/DO 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2679 GND 17_9/a_26_538# 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2680 17_9/DATA 17_9/a_420_786# 17_9/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2681 17_9/DIB 17_9/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2682 17_9/a_62_902# 17_9/a_26_538# 17_9/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2683 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2684 17_9/DI 17_9/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2685 Vdd 17_9/DO 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2686 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2687 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2688 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2689 Vdd 17_9/a_58_538# 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2690 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2691 GND 17_9/a_26_538# 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2692 17_9/a_62_902# 17_9/a_58_538# 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2693 17_9/DIB 17_9/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2694 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2695 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2696 17_9/a_62_82# 17_9/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2697 17_9/DI 17_9/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2698 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2699 17_9/a_62_82# 17_9/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2700 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2701 17_9/DATA 17_9/a_252_786# 17_9/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2702 Vdd 17_9/a_58_538# 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2703 17_9/a_62_82# 17_9/a_26_538# 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2704 GND 17_9/DATA 17_9/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2705 GND 17_9/DIB 17_9/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2706 17_9/a_62_902# 17_9/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2707 17_9/a_62_902# 17_9/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2708 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2709 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2710 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2711 17_9/a_62_82# 17_9/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2712 17_9/a_62_82# 17_9/a_58_538# 17_9/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2713 Vdd 17_9/DATA 17_9/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2714 Vdd 17_9/DIB 17_9/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2715 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2716 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2717 17_9/a_62_902# 17_9/a_26_538# 17_9/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2718 17_9/DIB 17_9/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2719 17_9/DI 17_9/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2720 17_9/a_62_902# 17_9/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2721 GND 17_9/DO 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2722 GND 17_9/DO 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2723 17_9/a_58_538# 17_9/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2724 17_9/a_62_902# 17_9/a_58_538# 17_9/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2725 17_9/DI 17_9/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2726 Vdd 17_9/DO 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2727 17_9/DIB 17_9/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2728 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2729 17_9/DIB 17_9/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2730 17_9/DI 17_9/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2731 GND 17_9/DATA 17_9/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2732 17_9/a_58_538# 17_9/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2733 Vdd 17_9/DO 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2734 17_9/a_62_82# 17_9/a_26_538# 17_9/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2735 GND 17_9/DIB 17_9/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2736 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2737 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2738 17_9/DIB 17_9/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2739 17_9/DI 17_9/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2740 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2741 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2742 17_9/a_62_82# 17_9/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2743 GND 17_9/a_62_82# 17_9/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2744 GND 17_9/OEN 17_9/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2745 17_9/a_62_82# 17_9/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2746 Vdd 17_9/DATA 17_9/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2747 Vdd 17_9/DIB 17_9/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2748 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2749 17_9/DATA 17_9/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2750 Vdd 17_9/a_62_902# 17_9/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2751 GND 17_9/DATA 17_9/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2752 GND 17_9/DIB 17_9/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2753 17_9/a_62_902# 17_9/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2754 Vdd 17_9/OEN 17_9/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2755 17_9/a_62_902# 17_9/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2756 17_9/a_62_82# 17_9/a_58_538# 17_9/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2757 Vdd 17_9/DATA 17_9/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2758 Vdd 17_9/DIB 17_9/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2759 17_9/DATA 17_9/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2760 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.4n ps=0.284m
M2761 Vdd GND GND GND nfet w=200 l=6
+  ad=8.4n pd=0.284m as=3.6n ps=0.236m
M2762 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M2763 Vdd GND GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M2764 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.436m as=8.4n ps=0.284m
M2765 Vdd GND GND GND nfet w=200 l=6
+  ad=8.4n pd=0.284m as=3.6n ps=0.236m
M2766 Vdd GND GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M2767 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M2768 Vdd GND GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.236m
M2769 Vdd GND GND GND nfet w=200 l=6
+  ad=8.2n pd=0.282m as=3.6n ps=0.436m
M2770 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M2771 GND GND Vdd GND nfet w=200 l=6
+  ad=3.6n pd=0.236m as=8.2n ps=0.282m
M2772 GND 17_30/DO 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2773 GND 17_30/a_26_538# 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2774 17_30/DATA 17_30/a_420_786# 17_30/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2775 17_30/DIB 17_30/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2776 17_30/a_62_902# 17_30/a_26_538# 17_30/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2777 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2778 17_30/DI 17_30/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2779 Vdd 17_30/DO 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2780 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2781 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2782 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2783 Vdd 17_30/a_58_538# 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2784 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2785 GND 17_30/a_26_538# 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2786 17_30/a_62_902# 17_30/a_58_538# 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2787 17_30/DIB 17_30/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2788 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2789 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2790 17_30/a_62_82# 17_30/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2791 17_30/DI 17_30/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2792 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2793 17_30/a_62_82# 17_30/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2794 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2795 17_30/DATA 17_30/a_252_786# 17_30/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2796 Vdd 17_30/a_58_538# 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2797 17_30/a_62_82# 17_30/a_26_538# 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2798 GND 17_30/DATA 17_30/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2799 GND 17_30/DIB 17_30/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2800 17_30/a_62_902# 17_30/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2801 17_30/a_62_902# 17_30/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2802 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2803 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2804 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2805 17_30/a_62_82# 17_30/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2806 17_30/a_62_82# 17_30/a_58_538# 17_30/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2807 Vdd 17_30/DATA 17_30/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2808 Vdd 17_30/DIB 17_30/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2809 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2810 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2811 17_30/a_62_902# 17_30/a_26_538# 17_30/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2812 17_30/DIB 17_30/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2813 17_30/DI 17_30/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2814 17_30/a_62_902# 17_30/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2815 GND 17_30/DO 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2816 GND 17_30/DO 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2817 17_30/a_58_538# 17_30/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2818 17_30/a_62_902# 17_30/a_58_538# 17_30/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2819 17_30/DI 17_30/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2820 Vdd 17_30/DO 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2821 17_30/DIB 17_30/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2822 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2823 17_30/DIB 17_30/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2824 17_30/DI 17_30/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2825 GND 17_30/DATA 17_30/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2826 17_30/a_58_538# 17_30/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2827 Vdd 17_30/DO 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2828 17_30/a_62_82# 17_30/a_26_538# 17_30/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2829 GND 17_30/DIB 17_30/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2830 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2831 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2832 17_30/DIB 17_30/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2833 17_30/DI 17_30/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2834 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2835 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2836 17_30/a_62_82# 17_30/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2837 GND 17_30/a_62_82# 17_30/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2838 GND 17_30/OEN 17_30/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2839 17_30/a_62_82# 17_30/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2840 Vdd 17_30/DATA 17_30/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2841 Vdd 17_30/DIB 17_30/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2842 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2843 17_30/DATA 17_30/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2844 Vdd 17_30/a_62_902# 17_30/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2845 GND 17_30/DATA 17_30/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2846 GND 17_30/DIB 17_30/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2847 17_30/a_62_902# 17_30/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2848 Vdd 17_30/OEN 17_30/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2849 17_30/a_62_902# 17_30/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2850 17_30/a_62_82# 17_30/a_58_538# 17_30/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2851 Vdd 17_30/DATA 17_30/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2852 Vdd 17_30/DIB 17_30/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2853 17_30/DATA 17_30/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2854 GND 17_20/DO 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2855 GND 17_20/a_26_538# 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2856 17_20/DATA 17_20/a_420_786# 17_20/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2857 17_20/DIB 17_20/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2858 17_20/a_62_902# 17_20/a_26_538# 17_20/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2859 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2860 17_20/DI 17_20/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2861 Vdd 17_20/DO 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2862 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2863 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2864 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2865 Vdd 17_20/a_58_538# 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2866 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2867 GND 17_20/a_26_538# 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2868 17_20/a_62_902# 17_20/a_58_538# 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2869 17_20/DIB 17_20/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2870 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2871 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2872 17_20/a_62_82# 17_20/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2873 17_20/DI 17_20/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2874 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2875 17_20/a_62_82# 17_20/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2876 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2877 17_20/DATA 17_20/a_252_786# 17_20/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2878 Vdd 17_20/a_58_538# 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2879 17_20/a_62_82# 17_20/a_26_538# 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2880 GND 17_20/DATA 17_20/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2881 GND 17_20/DIB 17_20/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2882 17_20/a_62_902# 17_20/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2883 17_20/a_62_902# 17_20/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2884 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2885 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2886 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2887 17_20/a_62_82# 17_20/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2888 17_20/a_62_82# 17_20/a_58_538# 17_20/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2889 Vdd 17_20/DATA 17_20/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2890 Vdd 17_20/DIB 17_20/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2891 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2892 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2893 17_20/a_62_902# 17_20/a_26_538# 17_20/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2894 17_20/DIB 17_20/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2895 17_20/DI 17_20/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2896 17_20/a_62_902# 17_20/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2897 GND 17_20/DO 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2898 GND 17_20/DO 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2899 17_20/a_58_538# 17_20/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2900 17_20/a_62_902# 17_20/a_58_538# 17_20/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2901 17_20/DI 17_20/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2902 Vdd 17_20/DO 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2903 17_20/DIB 17_20/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2904 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2905 17_20/DIB 17_20/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2906 17_20/DI 17_20/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2907 GND 17_20/DATA 17_20/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2908 17_20/a_58_538# 17_20/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2909 Vdd 17_20/DO 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2910 17_20/a_62_82# 17_20/a_26_538# 17_20/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2911 GND 17_20/DIB 17_20/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2912 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2913 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2914 17_20/DIB 17_20/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2915 17_20/DI 17_20/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2916 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2917 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2918 17_20/a_62_82# 17_20/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2919 GND 17_20/a_62_82# 17_20/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2920 GND 17_20/OEN 17_20/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M2921 17_20/a_62_82# 17_20/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2922 Vdd 17_20/DATA 17_20/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2923 Vdd 17_20/DIB 17_20/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2924 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2925 17_20/DATA 17_20/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2926 Vdd 17_20/a_62_902# 17_20/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2927 GND 17_20/DATA 17_20/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2928 GND 17_20/DIB 17_20/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2929 17_20/a_62_902# 17_20/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2930 Vdd 17_20/OEN 17_20/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M2931 17_20/a_62_902# 17_20/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2932 17_20/a_62_82# 17_20/a_58_538# 17_20/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2933 Vdd 17_20/DATA 17_20/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2934 Vdd 17_20/DIB 17_20/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2935 17_20/DATA 17_20/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2936 GND 17_31/DO 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M2937 GND 17_31/a_26_538# 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2938 17_31/DATA 17_31/a_420_786# 17_31/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M2939 17_31/DIB 17_31/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2940 17_31/a_62_902# 17_31/a_26_538# 17_31/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M2941 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M2942 17_31/DI 17_31/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M2943 Vdd 17_31/DO 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2944 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M2945 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2946 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2947 Vdd 17_31/a_58_538# 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2948 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2949 GND 17_31/a_26_538# 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2950 17_31/a_62_902# 17_31/a_58_538# 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M2951 17_31/DIB 17_31/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2952 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2953 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2954 17_31/a_62_82# 17_31/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2955 17_31/DI 17_31/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M2956 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2957 17_31/a_62_82# 17_31/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2958 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2959 17_31/DATA 17_31/a_252_786# 17_31/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M2960 Vdd 17_31/a_58_538# 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2961 17_31/a_62_82# 17_31/a_26_538# 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2962 GND 17_31/DATA 17_31/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2963 GND 17_31/DIB 17_31/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2964 17_31/a_62_902# 17_31/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2965 17_31/a_62_902# 17_31/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2966 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2967 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2968 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2969 17_31/a_62_82# 17_31/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2970 17_31/a_62_82# 17_31/a_58_538# 17_31/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2971 Vdd 17_31/DATA 17_31/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2972 Vdd 17_31/DIB 17_31/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2973 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2974 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2975 17_31/a_62_902# 17_31/a_26_538# 17_31/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2976 17_31/DIB 17_31/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2977 17_31/DI 17_31/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2978 17_31/a_62_902# 17_31/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2979 GND 17_31/DO 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2980 GND 17_31/DO 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2981 17_31/a_58_538# 17_31/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M2982 17_31/a_62_902# 17_31/a_58_538# 17_31/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2983 17_31/DI 17_31/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2984 Vdd 17_31/DO 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2985 17_31/DIB 17_31/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2986 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2987 17_31/DIB 17_31/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2988 17_31/DI 17_31/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2989 GND 17_31/DATA 17_31/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2990 17_31/a_58_538# 17_31/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M2991 Vdd 17_31/DO 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2992 17_31/a_62_82# 17_31/a_26_538# 17_31/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2993 GND 17_31/DIB 17_31/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M2994 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2995 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2996 17_31/DIB 17_31/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2997 17_31/DI 17_31/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M2998 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M2999 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3000 17_31/a_62_82# 17_31/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3001 GND 17_31/a_62_82# 17_31/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3002 GND 17_31/OEN 17_31/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3003 17_31/a_62_82# 17_31/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3004 Vdd 17_31/DATA 17_31/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3005 Vdd 17_31/DIB 17_31/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3006 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3007 17_31/DATA 17_31/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3008 Vdd 17_31/a_62_902# 17_31/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3009 GND 17_31/DATA 17_31/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3010 GND 17_31/DIB 17_31/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3011 17_31/a_62_902# 17_31/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3012 Vdd 17_31/OEN 17_31/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3013 17_31/a_62_902# 17_31/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3014 17_31/a_62_82# 17_31/a_58_538# 17_31/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3015 Vdd 17_31/DATA 17_31/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3016 Vdd 17_31/DIB 17_31/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3017 17_31/DATA 17_31/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3018 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=6.799297u ps=0.39057
M3019 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3020 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3021 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3022 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3023 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3024 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3025 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3026 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3027 Vdd GND GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3028 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3029 GND GND Vdd GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3030 GND 17_10/DO 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3031 GND 17_10/a_26_538# 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3032 17_10/DATA 17_10/a_420_786# 17_10/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3033 17_10/DIB 17_10/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3034 17_10/a_62_902# 17_10/a_26_538# 17_10/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3035 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3036 17_10/DI 17_10/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3037 Vdd 17_10/DO 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3038 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3039 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3040 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3041 Vdd 17_10/a_58_538# 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3042 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3043 GND 17_10/a_26_538# 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3044 17_10/a_62_902# 17_10/a_58_538# 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3045 17_10/DIB 17_10/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3046 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3047 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3048 17_10/a_62_82# 17_10/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3049 17_10/DI 17_10/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3050 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3051 17_10/a_62_82# 17_10/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3052 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3053 17_10/DATA 17_10/a_252_786# 17_10/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3054 Vdd 17_10/a_58_538# 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3055 17_10/a_62_82# 17_10/a_26_538# 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3056 GND 17_10/DATA 17_10/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3057 GND 17_10/DIB 17_10/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3058 17_10/a_62_902# 17_10/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3059 17_10/a_62_902# 17_10/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3060 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3061 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3062 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3063 17_10/a_62_82# 17_10/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3064 17_10/a_62_82# 17_10/a_58_538# 17_10/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3065 Vdd 17_10/DATA 17_10/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3066 Vdd 17_10/DIB 17_10/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3067 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3068 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3069 17_10/a_62_902# 17_10/a_26_538# 17_10/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3070 17_10/DIB 17_10/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3071 17_10/DI 17_10/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3072 17_10/a_62_902# 17_10/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3073 GND 17_10/DO 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3074 GND 17_10/DO 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3075 17_10/a_58_538# 17_10/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3076 17_10/a_62_902# 17_10/a_58_538# 17_10/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3077 17_10/DI 17_10/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3078 Vdd 17_10/DO 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3079 17_10/DIB 17_10/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3080 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3081 17_10/DIB 17_10/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3082 17_10/DI 17_10/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3083 GND 17_10/DATA 17_10/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3084 17_10/a_58_538# 17_10/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3085 Vdd 17_10/DO 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3086 17_10/a_62_82# 17_10/a_26_538# 17_10/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3087 GND 17_10/DIB 17_10/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3088 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3089 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3090 17_10/DIB 17_10/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3091 17_10/DI 17_10/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3092 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3093 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3094 17_10/a_62_82# 17_10/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3095 GND 17_10/a_62_82# 17_10/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3096 GND 17_10/OEN 17_10/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3097 17_10/a_62_82# 17_10/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3098 Vdd 17_10/DATA 17_10/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3099 Vdd 17_10/DIB 17_10/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3100 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3101 17_10/DATA 17_10/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3102 Vdd 17_10/a_62_902# 17_10/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3103 GND 17_10/DATA 17_10/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3104 GND 17_10/DIB 17_10/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3105 17_10/a_62_902# 17_10/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3106 Vdd 17_10/OEN 17_10/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3107 17_10/a_62_902# 17_10/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3108 17_10/a_62_82# 17_10/a_58_538# 17_10/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3109 Vdd 17_10/DATA 17_10/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3110 Vdd 17_10/DIB 17_10/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3111 17_10/DATA 17_10/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3112 GND 17_21/DO 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3113 GND 17_21/a_26_538# 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3114 17_21/DATA 17_21/a_420_786# 17_21/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3115 17_21/DIB 17_21/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3116 17_21/a_62_902# 17_21/a_26_538# 17_21/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3117 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3118 17_21/DI 17_21/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3119 Vdd 17_21/DO 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3120 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3121 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3122 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3123 Vdd 17_21/a_58_538# 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3124 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3125 GND 17_21/a_26_538# 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3126 17_21/a_62_902# 17_21/a_58_538# 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3127 17_21/DIB 17_21/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3128 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3129 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3130 17_21/a_62_82# 17_21/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3131 17_21/DI 17_21/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3132 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3133 17_21/a_62_82# 17_21/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3134 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3135 17_21/DATA 17_21/a_252_786# 17_21/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3136 Vdd 17_21/a_58_538# 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3137 17_21/a_62_82# 17_21/a_26_538# 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3138 GND 17_21/DATA 17_21/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3139 GND 17_21/DIB 17_21/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3140 17_21/a_62_902# 17_21/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3141 17_21/a_62_902# 17_21/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3142 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3143 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3144 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3145 17_21/a_62_82# 17_21/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3146 17_21/a_62_82# 17_21/a_58_538# 17_21/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3147 Vdd 17_21/DATA 17_21/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3148 Vdd 17_21/DIB 17_21/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3149 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3150 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3151 17_21/a_62_902# 17_21/a_26_538# 17_21/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3152 17_21/DIB 17_21/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3153 17_21/DI 17_21/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3154 17_21/a_62_902# 17_21/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3155 GND 17_21/DO 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3156 GND 17_21/DO 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3157 17_21/a_58_538# 17_21/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3158 17_21/a_62_902# 17_21/a_58_538# 17_21/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3159 17_21/DI 17_21/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3160 Vdd 17_21/DO 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3161 17_21/DIB 17_21/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3162 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3163 17_21/DIB 17_21/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3164 17_21/DI 17_21/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3165 GND 17_21/DATA 17_21/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3166 17_21/a_58_538# 17_21/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3167 Vdd 17_21/DO 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3168 17_21/a_62_82# 17_21/a_26_538# 17_21/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3169 GND 17_21/DIB 17_21/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3170 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3171 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3172 17_21/DIB 17_21/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3173 17_21/DI 17_21/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3174 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3175 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3176 17_21/a_62_82# 17_21/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3177 GND 17_21/a_62_82# 17_21/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3178 GND 17_21/OEN 17_21/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3179 17_21/a_62_82# 17_21/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3180 Vdd 17_21/DATA 17_21/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3181 Vdd 17_21/DIB 17_21/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3182 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3183 17_21/DATA 17_21/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3184 Vdd 17_21/a_62_902# 17_21/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3185 GND 17_21/DATA 17_21/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3186 GND 17_21/DIB 17_21/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3187 17_21/a_62_902# 17_21/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3188 Vdd 17_21/OEN 17_21/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3189 17_21/a_62_902# 17_21/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3190 17_21/a_62_82# 17_21/a_58_538# 17_21/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3191 Vdd 17_21/DATA 17_21/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3192 Vdd 17_21/DIB 17_21/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3193 17_21/DATA 17_21/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3194 GND 17_32/DO 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3195 GND 17_32/a_26_538# 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3196 17_32/DATA 17_32/a_420_786# 17_32/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3197 17_32/DIB 17_32/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3198 17_32/a_62_902# 17_32/a_26_538# 17_32/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3199 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3200 17_32/DI 17_32/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3201 Vdd 17_32/DO 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3202 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3203 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3204 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3205 Vdd 17_32/a_58_538# 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3206 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3207 GND 17_32/a_26_538# 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3208 17_32/a_62_902# 17_32/a_58_538# 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3209 17_32/DIB 17_32/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3210 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3211 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3212 17_32/a_62_82# 17_32/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3213 17_32/DI 17_32/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3214 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3215 17_32/a_62_82# 17_32/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3216 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3217 17_32/DATA 17_32/a_252_786# 17_32/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3218 Vdd 17_32/a_58_538# 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3219 17_32/a_62_82# 17_32/a_26_538# 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3220 GND 17_32/DATA 17_32/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3221 GND 17_32/DIB 17_32/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3222 17_32/a_62_902# 17_32/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3223 17_32/a_62_902# 17_32/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3224 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3225 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3226 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3227 17_32/a_62_82# 17_32/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3228 17_32/a_62_82# 17_32/a_58_538# 17_32/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3229 Vdd 17_32/DATA 17_32/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3230 Vdd 17_32/DIB 17_32/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3231 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3232 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3233 17_32/a_62_902# 17_32/a_26_538# 17_32/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3234 17_32/DIB 17_32/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3235 17_32/DI 17_32/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3236 17_32/a_62_902# 17_32/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3237 GND 17_32/DO 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3238 GND 17_32/DO 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3239 17_32/a_58_538# 17_32/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3240 17_32/a_62_902# 17_32/a_58_538# 17_32/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3241 17_32/DI 17_32/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3242 Vdd 17_32/DO 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3243 17_32/DIB 17_32/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3244 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3245 17_32/DIB 17_32/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3246 17_32/DI 17_32/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3247 GND 17_32/DATA 17_32/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3248 17_32/a_58_538# 17_32/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3249 Vdd 17_32/DO 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3250 17_32/a_62_82# 17_32/a_26_538# 17_32/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3251 GND 17_32/DIB 17_32/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3252 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3253 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3254 17_32/DIB 17_32/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3255 17_32/DI 17_32/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3256 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3257 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3258 17_32/a_62_82# 17_32/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3259 GND 17_32/a_62_82# 17_32/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3260 GND 17_32/OEN 17_32/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3261 17_32/a_62_82# 17_32/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3262 Vdd 17_32/DATA 17_32/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3263 Vdd 17_32/DIB 17_32/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3264 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3265 17_32/DATA 17_32/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3266 Vdd 17_32/a_62_902# 17_32/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3267 GND 17_32/DATA 17_32/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3268 GND 17_32/DIB 17_32/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3269 17_32/a_62_902# 17_32/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3270 Vdd 17_32/OEN 17_32/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3271 17_32/a_62_902# 17_32/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3272 17_32/a_62_82# 17_32/a_58_538# 17_32/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3273 Vdd 17_32/DATA 17_32/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3274 Vdd 17_32/DIB 17_32/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3275 17_32/DATA 17_32/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3276 GND 17_11/DO 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3277 GND 17_11/a_26_538# 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3278 17_11/DATA 17_11/a_420_786# 17_11/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3279 17_11/DIB 17_11/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3280 17_11/a_62_902# 17_11/a_26_538# 17_11/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3281 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3282 17_11/DI 17_11/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3283 Vdd 17_11/DO 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3284 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3285 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3286 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3287 Vdd 17_11/a_58_538# 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3288 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3289 GND 17_11/a_26_538# 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3290 17_11/a_62_902# 17_11/a_58_538# 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3291 17_11/DIB 17_11/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3292 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3293 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3294 17_11/a_62_82# 17_11/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3295 17_11/DI 17_11/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3296 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3297 17_11/a_62_82# 17_11/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3298 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3299 17_11/DATA 17_11/a_252_786# 17_11/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3300 Vdd 17_11/a_58_538# 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3301 17_11/a_62_82# 17_11/a_26_538# 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3302 GND 17_11/DATA 17_11/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3303 GND 17_11/DIB 17_11/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3304 17_11/a_62_902# 17_11/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3305 17_11/a_62_902# 17_11/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3306 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3307 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3308 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3309 17_11/a_62_82# 17_11/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3310 17_11/a_62_82# 17_11/a_58_538# 17_11/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3311 Vdd 17_11/DATA 17_11/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3312 Vdd 17_11/DIB 17_11/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3313 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3314 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3315 17_11/a_62_902# 17_11/a_26_538# 17_11/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3316 17_11/DIB 17_11/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3317 17_11/DI 17_11/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3318 17_11/a_62_902# 17_11/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3319 GND 17_11/DO 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3320 GND 17_11/DO 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3321 17_11/a_58_538# 17_11/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3322 17_11/a_62_902# 17_11/a_58_538# 17_11/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3323 17_11/DI 17_11/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3324 Vdd 17_11/DO 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3325 17_11/DIB 17_11/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3326 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3327 17_11/DIB 17_11/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3328 17_11/DI 17_11/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3329 GND 17_11/DATA 17_11/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3330 17_11/a_58_538# 17_11/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3331 Vdd 17_11/DO 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3332 17_11/a_62_82# 17_11/a_26_538# 17_11/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3333 GND 17_11/DIB 17_11/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3334 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3335 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3336 17_11/DIB 17_11/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3337 17_11/DI 17_11/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3338 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3339 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3340 17_11/a_62_82# 17_11/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3341 GND 17_11/a_62_82# 17_11/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3342 GND 17_11/OEN 17_11/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3343 17_11/a_62_82# 17_11/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3344 Vdd 17_11/DATA 17_11/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3345 Vdd 17_11/DIB 17_11/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3346 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3347 17_11/DATA 17_11/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3348 Vdd 17_11/a_62_902# 17_11/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3349 GND 17_11/DATA 17_11/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3350 GND 17_11/DIB 17_11/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3351 17_11/a_62_902# 17_11/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3352 Vdd 17_11/OEN 17_11/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3353 17_11/a_62_902# 17_11/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3354 17_11/a_62_82# 17_11/a_58_538# 17_11/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3355 Vdd 17_11/DATA 17_11/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3356 Vdd 17_11/DIB 17_11/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3357 17_11/DATA 17_11/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3358 GND 17_22/DO 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3359 GND 17_22/a_26_538# 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3360 17_22/DATA 17_22/a_420_786# 17_22/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3361 17_22/DIB 17_22/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3362 17_22/a_62_902# 17_22/a_26_538# 17_22/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3363 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3364 17_22/DI 17_22/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3365 Vdd 17_22/DO 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3366 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3367 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3368 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3369 Vdd 17_22/a_58_538# 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3370 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3371 GND 17_22/a_26_538# 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3372 17_22/a_62_902# 17_22/a_58_538# 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3373 17_22/DIB 17_22/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3374 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3375 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3376 17_22/a_62_82# 17_22/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3377 17_22/DI 17_22/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3378 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3379 17_22/a_62_82# 17_22/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3380 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3381 17_22/DATA 17_22/a_252_786# 17_22/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3382 Vdd 17_22/a_58_538# 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3383 17_22/a_62_82# 17_22/a_26_538# 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3384 GND 17_22/DATA 17_22/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3385 GND 17_22/DIB 17_22/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3386 17_22/a_62_902# 17_22/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3387 17_22/a_62_902# 17_22/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3388 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3389 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3390 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3391 17_22/a_62_82# 17_22/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3392 17_22/a_62_82# 17_22/a_58_538# 17_22/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3393 Vdd 17_22/DATA 17_22/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3394 Vdd 17_22/DIB 17_22/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3395 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3396 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3397 17_22/a_62_902# 17_22/a_26_538# 17_22/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3398 17_22/DIB 17_22/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3399 17_22/DI 17_22/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3400 17_22/a_62_902# 17_22/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3401 GND 17_22/DO 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3402 GND 17_22/DO 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3403 17_22/a_58_538# 17_22/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3404 17_22/a_62_902# 17_22/a_58_538# 17_22/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3405 17_22/DI 17_22/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3406 Vdd 17_22/DO 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3407 17_22/DIB 17_22/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3408 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3409 17_22/DIB 17_22/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3410 17_22/DI 17_22/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3411 GND 17_22/DATA 17_22/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3412 17_22/a_58_538# 17_22/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3413 Vdd 17_22/DO 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3414 17_22/a_62_82# 17_22/a_26_538# 17_22/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3415 GND 17_22/DIB 17_22/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3416 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3417 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3418 17_22/DIB 17_22/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3419 17_22/DI 17_22/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3420 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3421 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3422 17_22/a_62_82# 17_22/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3423 GND 17_22/a_62_82# 17_22/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3424 GND 17_22/OEN 17_22/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3425 17_22/a_62_82# 17_22/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3426 Vdd 17_22/DATA 17_22/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3427 Vdd 17_22/DIB 17_22/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3428 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3429 17_22/DATA 17_22/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3430 Vdd 17_22/a_62_902# 17_22/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3431 GND 17_22/DATA 17_22/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3432 GND 17_22/DIB 17_22/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3433 17_22/a_62_902# 17_22/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3434 Vdd 17_22/OEN 17_22/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3435 17_22/a_62_902# 17_22/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3436 17_22/a_62_82# 17_22/a_58_538# 17_22/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3437 Vdd 17_22/DATA 17_22/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3438 Vdd 17_22/DIB 17_22/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3439 17_22/DATA 17_22/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3440 GND 17_33/DO 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3441 GND 17_33/a_26_538# 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3442 17_33/DATA 17_33/a_420_786# 17_33/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3443 17_33/DIB 17_33/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3444 17_33/a_62_902# 17_33/a_26_538# 17_33/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3445 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3446 17_33/DI 17_33/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3447 Vdd 17_33/DO 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3448 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3449 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3450 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3451 Vdd 17_33/a_58_538# 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3452 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3453 GND 17_33/a_26_538# 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3454 17_33/a_62_902# 17_33/a_58_538# 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3455 17_33/DIB 17_33/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3456 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3457 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3458 17_33/a_62_82# 17_33/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3459 17_33/DI 17_33/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3460 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3461 17_33/a_62_82# 17_33/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3462 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3463 17_33/DATA 17_33/a_252_786# 17_33/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3464 Vdd 17_33/a_58_538# 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3465 17_33/a_62_82# 17_33/a_26_538# 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3466 GND 17_33/DATA 17_33/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3467 GND 17_33/DIB 17_33/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3468 17_33/a_62_902# 17_33/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3469 17_33/a_62_902# 17_33/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3470 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3471 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3472 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3473 17_33/a_62_82# 17_33/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3474 17_33/a_62_82# 17_33/a_58_538# 17_33/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3475 Vdd 17_33/DATA 17_33/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3476 Vdd 17_33/DIB 17_33/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3477 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3478 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3479 17_33/a_62_902# 17_33/a_26_538# 17_33/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3480 17_33/DIB 17_33/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3481 17_33/DI 17_33/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3482 17_33/a_62_902# 17_33/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3483 GND 17_33/DO 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3484 GND 17_33/DO 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3485 17_33/a_58_538# 17_33/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3486 17_33/a_62_902# 17_33/a_58_538# 17_33/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3487 17_33/DI 17_33/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3488 Vdd 17_33/DO 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3489 17_33/DIB 17_33/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3490 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3491 17_33/DIB 17_33/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3492 17_33/DI 17_33/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3493 GND 17_33/DATA 17_33/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3494 17_33/a_58_538# 17_33/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3495 Vdd 17_33/DO 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3496 17_33/a_62_82# 17_33/a_26_538# 17_33/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3497 GND 17_33/DIB 17_33/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3498 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3499 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3500 17_33/DIB 17_33/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3501 17_33/DI 17_33/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3502 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3503 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3504 17_33/a_62_82# 17_33/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3505 GND 17_33/a_62_82# 17_33/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3506 GND 17_33/OEN 17_33/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3507 17_33/a_62_82# 17_33/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3508 Vdd 17_33/DATA 17_33/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3509 Vdd 17_33/DIB 17_33/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3510 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3511 17_33/DATA 17_33/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3512 Vdd 17_33/a_62_902# 17_33/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3513 GND 17_33/DATA 17_33/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3514 GND 17_33/DIB 17_33/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3515 17_33/a_62_902# 17_33/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3516 Vdd 17_33/OEN 17_33/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3517 17_33/a_62_902# 17_33/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3518 17_33/a_62_82# 17_33/a_58_538# 17_33/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3519 Vdd 17_33/DATA 17_33/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3520 Vdd 17_33/DIB 17_33/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3521 17_33/DATA 17_33/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3522 GND 17_12/DO 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3523 GND 17_12/a_26_538# 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3524 17_12/DATA 17_12/a_420_786# 17_12/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3525 17_12/DIB 17_12/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3526 17_12/a_62_902# 17_12/a_26_538# 17_12/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3527 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3528 17_12/DI 17_12/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3529 Vdd 17_12/DO 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3530 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3531 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3532 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3533 Vdd 17_12/a_58_538# 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3534 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3535 GND 17_12/a_26_538# 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3536 17_12/a_62_902# 17_12/a_58_538# 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3537 17_12/DIB 17_12/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3538 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3539 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3540 17_12/a_62_82# 17_12/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3541 17_12/DI 17_12/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3542 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3543 17_12/a_62_82# 17_12/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3544 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3545 17_12/DATA 17_12/a_252_786# 17_12/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3546 Vdd 17_12/a_58_538# 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3547 17_12/a_62_82# 17_12/a_26_538# 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3548 GND 17_12/DATA 17_12/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3549 GND 17_12/DIB 17_12/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3550 17_12/a_62_902# 17_12/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3551 17_12/a_62_902# 17_12/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3552 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3553 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3554 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3555 17_12/a_62_82# 17_12/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3556 17_12/a_62_82# 17_12/a_58_538# 17_12/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3557 Vdd 17_12/DATA 17_12/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3558 Vdd 17_12/DIB 17_12/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3559 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3560 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3561 17_12/a_62_902# 17_12/a_26_538# 17_12/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3562 17_12/DIB 17_12/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3563 17_12/DI 17_12/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3564 17_12/a_62_902# 17_12/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3565 GND 17_12/DO 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3566 GND 17_12/DO 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3567 17_12/a_58_538# 17_12/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3568 17_12/a_62_902# 17_12/a_58_538# 17_12/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3569 17_12/DI 17_12/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3570 Vdd 17_12/DO 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3571 17_12/DIB 17_12/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3572 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3573 17_12/DIB 17_12/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3574 17_12/DI 17_12/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3575 GND 17_12/DATA 17_12/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3576 17_12/a_58_538# 17_12/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3577 Vdd 17_12/DO 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3578 17_12/a_62_82# 17_12/a_26_538# 17_12/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3579 GND 17_12/DIB 17_12/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3580 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3581 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3582 17_12/DIB 17_12/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3583 17_12/DI 17_12/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3584 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3585 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3586 17_12/a_62_82# 17_12/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3587 GND 17_12/a_62_82# 17_12/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3588 GND 17_12/OEN 17_12/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3589 17_12/a_62_82# 17_12/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3590 Vdd 17_12/DATA 17_12/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3591 Vdd 17_12/DIB 17_12/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3592 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3593 17_12/DATA 17_12/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3594 Vdd 17_12/a_62_902# 17_12/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3595 GND 17_12/DATA 17_12/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3596 GND 17_12/DIB 17_12/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3597 17_12/a_62_902# 17_12/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3598 Vdd 17_12/OEN 17_12/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3599 17_12/a_62_902# 17_12/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3600 17_12/a_62_82# 17_12/a_58_538# 17_12/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3601 Vdd 17_12/DATA 17_12/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3602 Vdd 17_12/DIB 17_12/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3603 17_12/DATA 17_12/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3604 GND 17_13/DO 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3605 GND 17_13/a_26_538# 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3606 17_13/DATA 17_13/a_420_786# 17_13/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3607 17_13/DIB 17_13/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3608 17_13/a_62_902# 17_13/a_26_538# 17_13/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3609 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3610 17_13/DI 17_13/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3611 Vdd 17_13/DO 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3612 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3613 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3614 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3615 Vdd 17_13/a_58_538# 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3616 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3617 GND 17_13/a_26_538# 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3618 17_13/a_62_902# 17_13/a_58_538# 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3619 17_13/DIB 17_13/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3620 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3621 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3622 17_13/a_62_82# 17_13/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3623 17_13/DI 17_13/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3624 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3625 17_13/a_62_82# 17_13/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3626 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3627 17_13/DATA 17_13/a_252_786# 17_13/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3628 Vdd 17_13/a_58_538# 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3629 17_13/a_62_82# 17_13/a_26_538# 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3630 GND 17_13/DATA 17_13/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3631 GND 17_13/DIB 17_13/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3632 17_13/a_62_902# 17_13/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3633 17_13/a_62_902# 17_13/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3634 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3635 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3636 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3637 17_13/a_62_82# 17_13/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3638 17_13/a_62_82# 17_13/a_58_538# 17_13/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3639 Vdd 17_13/DATA 17_13/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3640 Vdd 17_13/DIB 17_13/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3641 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3642 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3643 17_13/a_62_902# 17_13/a_26_538# 17_13/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3644 17_13/DIB 17_13/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3645 17_13/DI 17_13/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3646 17_13/a_62_902# 17_13/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3647 GND 17_13/DO 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3648 GND 17_13/DO 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3649 17_13/a_58_538# 17_13/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3650 17_13/a_62_902# 17_13/a_58_538# 17_13/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3651 17_13/DI 17_13/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3652 Vdd 17_13/DO 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3653 17_13/DIB 17_13/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3654 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3655 17_13/DIB 17_13/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3656 17_13/DI 17_13/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3657 GND 17_13/DATA 17_13/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3658 17_13/a_58_538# 17_13/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3659 Vdd 17_13/DO 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3660 17_13/a_62_82# 17_13/a_26_538# 17_13/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3661 GND 17_13/DIB 17_13/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3662 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3663 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3664 17_13/DIB 17_13/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3665 17_13/DI 17_13/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3666 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3667 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3668 17_13/a_62_82# 17_13/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3669 GND 17_13/a_62_82# 17_13/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3670 GND 17_13/OEN 17_13/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3671 17_13/a_62_82# 17_13/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3672 Vdd 17_13/DATA 17_13/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3673 Vdd 17_13/DIB 17_13/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3674 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3675 17_13/DATA 17_13/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3676 Vdd 17_13/a_62_902# 17_13/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3677 GND 17_13/DATA 17_13/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3678 GND 17_13/DIB 17_13/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3679 17_13/a_62_902# 17_13/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3680 Vdd 17_13/OEN 17_13/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3681 17_13/a_62_902# 17_13/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3682 17_13/a_62_82# 17_13/a_58_538# 17_13/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3683 Vdd 17_13/DATA 17_13/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3684 Vdd 17_13/DIB 17_13/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3685 17_13/DATA 17_13/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3686 GND 17_23/DO 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3687 GND 17_23/a_26_538# 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3688 17_23/DATA 17_23/a_420_786# 17_23/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3689 17_23/DIB 17_23/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3690 17_23/a_62_902# 17_23/a_26_538# 17_23/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3691 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3692 17_23/DI 17_23/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3693 Vdd 17_23/DO 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3694 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3695 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3696 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3697 Vdd 17_23/a_58_538# 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3698 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3699 GND 17_23/a_26_538# 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3700 17_23/a_62_902# 17_23/a_58_538# 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3701 17_23/DIB 17_23/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3702 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3703 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3704 17_23/a_62_82# 17_23/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3705 17_23/DI 17_23/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3706 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3707 17_23/a_62_82# 17_23/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3708 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3709 17_23/DATA 17_23/a_252_786# 17_23/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3710 Vdd 17_23/a_58_538# 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3711 17_23/a_62_82# 17_23/a_26_538# 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3712 GND 17_23/DATA 17_23/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3713 GND 17_23/DIB 17_23/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3714 17_23/a_62_902# 17_23/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3715 17_23/a_62_902# 17_23/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3716 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3717 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3718 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3719 17_23/a_62_82# 17_23/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3720 17_23/a_62_82# 17_23/a_58_538# 17_23/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3721 Vdd 17_23/DATA 17_23/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3722 Vdd 17_23/DIB 17_23/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3723 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3724 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3725 17_23/a_62_902# 17_23/a_26_538# 17_23/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3726 17_23/DIB 17_23/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3727 17_23/DI 17_23/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3728 17_23/a_62_902# 17_23/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3729 GND 17_23/DO 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3730 GND 17_23/DO 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3731 17_23/a_58_538# 17_23/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3732 17_23/a_62_902# 17_23/a_58_538# 17_23/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3733 17_23/DI 17_23/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3734 Vdd 17_23/DO 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3735 17_23/DIB 17_23/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3736 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3737 17_23/DIB 17_23/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3738 17_23/DI 17_23/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3739 GND 17_23/DATA 17_23/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3740 17_23/a_58_538# 17_23/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3741 Vdd 17_23/DO 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3742 17_23/a_62_82# 17_23/a_26_538# 17_23/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3743 GND 17_23/DIB 17_23/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3744 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3745 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3746 17_23/DIB 17_23/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3747 17_23/DI 17_23/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3748 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3749 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3750 17_23/a_62_82# 17_23/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3751 GND 17_23/a_62_82# 17_23/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3752 GND 17_23/OEN 17_23/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3753 17_23/a_62_82# 17_23/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3754 Vdd 17_23/DATA 17_23/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3755 Vdd 17_23/DIB 17_23/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3756 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3757 17_23/DATA 17_23/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3758 Vdd 17_23/a_62_902# 17_23/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3759 GND 17_23/DATA 17_23/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3760 GND 17_23/DIB 17_23/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3761 17_23/a_62_902# 17_23/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3762 Vdd 17_23/OEN 17_23/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3763 17_23/a_62_902# 17_23/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3764 17_23/a_62_82# 17_23/a_58_538# 17_23/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3765 Vdd 17_23/DATA 17_23/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3766 Vdd 17_23/DIB 17_23/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3767 17_23/DATA 17_23/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3768 GND 17_24/DO 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3769 GND 17_24/a_26_538# 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3770 17_24/DATA 17_24/a_420_786# 17_24/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3771 17_24/DIB 17_24/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3772 17_24/a_62_902# 17_24/a_26_538# 17_24/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3773 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3774 17_24/DI 17_24/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3775 Vdd 17_24/DO 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3776 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3777 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3778 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3779 Vdd 17_24/a_58_538# 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3780 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3781 GND 17_24/a_26_538# 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3782 17_24/a_62_902# 17_24/a_58_538# 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3783 17_24/DIB 17_24/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3784 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3785 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3786 17_24/a_62_82# 17_24/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3787 17_24/DI 17_24/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3788 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3789 17_24/a_62_82# 17_24/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3790 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3791 17_24/DATA 17_24/a_252_786# 17_24/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3792 Vdd 17_24/a_58_538# 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3793 17_24/a_62_82# 17_24/a_26_538# 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3794 GND 17_24/DATA 17_24/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3795 GND 17_24/DIB 17_24/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3796 17_24/a_62_902# 17_24/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3797 17_24/a_62_902# 17_24/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3798 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3799 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3800 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3801 17_24/a_62_82# 17_24/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3802 17_24/a_62_82# 17_24/a_58_538# 17_24/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3803 Vdd 17_24/DATA 17_24/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3804 Vdd 17_24/DIB 17_24/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3805 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3806 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3807 17_24/a_62_902# 17_24/a_26_538# 17_24/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3808 17_24/DIB 17_24/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3809 17_24/DI 17_24/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3810 17_24/a_62_902# 17_24/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3811 GND 17_24/DO 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3812 GND 17_24/DO 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3813 17_24/a_58_538# 17_24/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3814 17_24/a_62_902# 17_24/a_58_538# 17_24/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3815 17_24/DI 17_24/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3816 Vdd 17_24/DO 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3817 17_24/DIB 17_24/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3818 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3819 17_24/DIB 17_24/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3820 17_24/DI 17_24/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3821 GND 17_24/DATA 17_24/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3822 17_24/a_58_538# 17_24/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3823 Vdd 17_24/DO 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3824 17_24/a_62_82# 17_24/a_26_538# 17_24/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3825 GND 17_24/DIB 17_24/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3826 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3827 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3828 17_24/DIB 17_24/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3829 17_24/DI 17_24/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3830 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3831 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3832 17_24/a_62_82# 17_24/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3833 GND 17_24/a_62_82# 17_24/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3834 GND 17_24/OEN 17_24/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3835 17_24/a_62_82# 17_24/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3836 Vdd 17_24/DATA 17_24/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3837 Vdd 17_24/DIB 17_24/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3838 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3839 17_24/DATA 17_24/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3840 Vdd 17_24/a_62_902# 17_24/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3841 GND 17_24/DATA 17_24/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3842 GND 17_24/DIB 17_24/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3843 17_24/a_62_902# 17_24/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3844 Vdd 17_24/OEN 17_24/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3845 17_24/a_62_902# 17_24/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3846 17_24/a_62_82# 17_24/a_58_538# 17_24/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3847 Vdd 17_24/DATA 17_24/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3848 Vdd 17_24/DIB 17_24/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3849 17_24/DATA 17_24/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3850 GND 17_34/DO 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3851 GND 17_34/a_26_538# 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3852 17_34/DATA 17_34/a_420_786# 17_34/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3853 17_34/DIB 17_34/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3854 17_34/a_62_902# 17_34/a_26_538# 17_34/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3855 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3856 17_34/DI 17_34/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3857 Vdd 17_34/DO 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3858 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3859 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3860 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3861 Vdd 17_34/a_58_538# 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3862 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3863 GND 17_34/a_26_538# 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3864 17_34/a_62_902# 17_34/a_58_538# 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3865 17_34/DIB 17_34/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3866 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3867 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3868 17_34/a_62_82# 17_34/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3869 17_34/DI 17_34/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3870 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3871 17_34/a_62_82# 17_34/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3872 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3873 17_34/DATA 17_34/a_252_786# 17_34/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3874 Vdd 17_34/a_58_538# 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3875 17_34/a_62_82# 17_34/a_26_538# 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3876 GND 17_34/DATA 17_34/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3877 GND 17_34/DIB 17_34/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3878 17_34/a_62_902# 17_34/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3879 17_34/a_62_902# 17_34/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3880 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3881 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3882 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3883 17_34/a_62_82# 17_34/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3884 17_34/a_62_82# 17_34/a_58_538# 17_34/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3885 Vdd 17_34/DATA 17_34/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3886 Vdd 17_34/DIB 17_34/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3887 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3888 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3889 17_34/a_62_902# 17_34/a_26_538# 17_34/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3890 17_34/DIB 17_34/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3891 17_34/DI 17_34/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3892 17_34/a_62_902# 17_34/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3893 GND 17_34/DO 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3894 GND 17_34/DO 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3895 17_34/a_58_538# 17_34/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3896 17_34/a_62_902# 17_34/a_58_538# 17_34/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3897 17_34/DI 17_34/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3898 Vdd 17_34/DO 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3899 17_34/DIB 17_34/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3900 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3901 17_34/DIB 17_34/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3902 17_34/DI 17_34/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3903 GND 17_34/DATA 17_34/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3904 17_34/a_58_538# 17_34/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3905 Vdd 17_34/DO 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3906 17_34/a_62_82# 17_34/a_26_538# 17_34/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3907 GND 17_34/DIB 17_34/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3908 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3909 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3910 17_34/DIB 17_34/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3911 17_34/DI 17_34/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3912 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3913 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3914 17_34/a_62_82# 17_34/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3915 GND 17_34/a_62_82# 17_34/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3916 GND 17_34/OEN 17_34/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3917 17_34/a_62_82# 17_34/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3918 Vdd 17_34/DATA 17_34/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3919 Vdd 17_34/DIB 17_34/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3920 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3921 17_34/DATA 17_34/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3922 Vdd 17_34/a_62_902# 17_34/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3923 GND 17_34/DATA 17_34/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3924 GND 17_34/DIB 17_34/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3925 17_34/a_62_902# 17_34/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3926 Vdd 17_34/OEN 17_34/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M3927 17_34/a_62_902# 17_34/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3928 17_34/a_62_82# 17_34/a_58_538# 17_34/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3929 Vdd 17_34/DATA 17_34/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3930 Vdd 17_34/DIB 17_34/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3931 17_34/DATA 17_34/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3932 GND 17_35/DO 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=5.76n ps=1.152m
M3933 GND 17_35/a_26_538# 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3934 17_35/DATA 17_35/a_420_786# 17_35/DATA Gnd polyResistor w=20 l=128
+  ad=7.7n pd=2.824m as=0 ps=0
M3935 17_35/DIB 17_35/DATA GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3936 17_35/a_62_902# 17_35/a_26_538# 17_35/a_62_82# Vdd pfet w=104 l=4
+  ad=9.984n pd=1.856m as=2.496n ps=0.464m
M3937 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=97.6n ps=3.376m
M3938 17_35/DI 17_35/DIB GND Gnd nfet w=60 l=4
+  ad=2.16n pd=0.432m as=0 ps=0
M3939 Vdd 17_35/DO 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3940 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=99.200005n ps=3.392m
M3941 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3942 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3943 Vdd 17_35/a_58_538# 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3944 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3945 GND 17_35/a_26_538# 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3946 17_35/a_62_902# 17_35/a_58_538# 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=1.44n pd=0.288m as=0 ps=0
M3947 17_35/DIB 17_35/DATA Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3948 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3949 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3950 17_35/a_62_82# 17_35/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3951 17_35/DI 17_35/DIB Vdd Vdd pfet w=104 l=4
+  ad=3.744n pd=0.696m as=0 ps=0
M3952 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3953 17_35/a_62_82# 17_35/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3954 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3955 17_35/DATA 17_35/a_252_786# 17_35/DATA Gnd polyResistor w=20 l=130
+  ad=0 pd=0 as=0 ps=0
M3956 Vdd 17_35/a_58_538# 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3957 17_35/a_62_82# 17_35/a_26_538# 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3958 GND 17_35/DATA 17_35/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3959 GND 17_35/DIB 17_35/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3960 17_35/a_62_902# 17_35/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3961 17_35/a_62_902# 17_35/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3962 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3963 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3964 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3965 17_35/a_62_82# 17_35/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3966 17_35/a_62_82# 17_35/a_58_538# 17_35/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3967 Vdd 17_35/DATA 17_35/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3968 Vdd 17_35/DIB 17_35/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3969 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3970 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3971 17_35/a_62_902# 17_35/a_26_538# 17_35/a_62_82# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3972 17_35/DIB 17_35/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3973 17_35/DI 17_35/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3974 17_35/a_62_902# 17_35/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3975 GND 17_35/DO 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3976 GND 17_35/DO 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3977 17_35/a_58_538# 17_35/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0.72n pd=0.144m as=0 ps=0
M3978 17_35/a_62_902# 17_35/a_58_538# 17_35/a_62_82# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3979 17_35/DI 17_35/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3980 Vdd 17_35/DO 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3981 17_35/DIB 17_35/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3982 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3983 17_35/DIB 17_35/DATA GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3984 17_35/DI 17_35/DIB GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3985 GND 17_35/DATA 17_35/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3986 17_35/a_58_538# 17_35/a_26_538# Vdd Vdd pfet w=104 l=4
+  ad=1.248n pd=0.232m as=0 ps=0
M3987 Vdd 17_35/DO 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3988 17_35/a_62_82# 17_35/a_26_538# 17_35/a_62_902# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3989 GND 17_35/DIB 17_35/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3990 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3991 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3992 17_35/DIB 17_35/DATA Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3993 17_35/DI 17_35/DIB Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M3994 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3995 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3996 17_35/a_62_82# 17_35/a_26_538# GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M3997 GND 17_35/a_62_82# 17_35/DATA GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M3998 GND 17_35/OEN 17_35/a_26_538# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0.72n ps=0.144m
M3999 17_35/a_62_82# 17_35/DO GND Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M4000 Vdd 17_35/DATA 17_35/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4001 Vdd 17_35/DIB 17_35/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4002 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M4003 17_35/DATA 17_35/a_62_902# Vdd Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M4004 Vdd 17_35/a_62_902# 17_35/DATA Vdd pfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
M4005 GND 17_35/DATA 17_35/DIB Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M4006 GND 17_35/DIB 17_35/DI Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M4007 17_35/a_62_902# 17_35/a_58_538# Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4008 Vdd 17_35/OEN 17_35/a_26_538# Vdd pfet w=104 l=4
+  ad=0 pd=0 as=1.248n ps=0.232m
M4009 17_35/a_62_902# 17_35/DO Vdd Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4010 17_35/a_62_82# 17_35/a_58_538# 17_35/a_62_902# Gnd nfet w=60 l=4
+  ad=0 pd=0 as=0 ps=0
M4011 Vdd 17_35/DATA 17_35/DIB Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4012 Vdd 17_35/DIB 17_35/DI Vdd pfet w=104 l=4
+  ad=0 pd=0 as=0 ps=0
M4013 17_35/DATA 17_35/a_62_82# GND GND nfet w=200 l=6
+  ad=0 pd=0 as=0 ps=0
C0 Vdd 17_26/DI 3.31488f
C1 GND 17_26/a_62_82# 48.660957f
C2 GND 17_24/OEN 4.46481f
C3 Vdd 17_24/DO 3.11769f
C4 17_5/a_420_786# p_d 2.95776f
C5 GND 17_33/DIB 6.35733f
C6 GND 17_21/m3_n72_n22# 32.78878f
C7 17_8/a_62_902# 17_8/DATA 6.99264f
C8 p_d 17_5/a_62_82# 8.056081f
C9 Vdd h 3.84291f
C10 17_26/a_62_902# 17_26/DATA 6.99264f
C11 Vdd 17_4/a_26_538# 3.76551f
C12 GND p_b 0.100362p
C13 17_12/a_252_786# 17_12/DATA 3.00456f
C14 GND 17_18/a_62_902# 2.79216f
C15 GND 17_10/a_26_538# 3.75903f
C16 GND 17_29/a_62_82# 48.660957f
C17 Vdd d 3.6576f
C18 GND 17_23/OEN 4.46481f
C19 Vdd 17_23/DO 3.11769f
C20 Vdd 17_18/DIB 6.39135f
C21 GND 17_18/a_58_538# 3.79746f
C22 GND 17_22/DIB 6.35733f
C23 GND 17_10/m3_n72_n22# 32.52166f
C24 17_14/a_26_538# Vdd 3.76551f
C25 17_14/DATA GND 0.100362p
C26 17_4/w_40_1480# p_b 66.6688f
C27 17_31/a_252_786# 17_31/DATA 3.00456f
C28 GND p_i 0.100362p
C29 Vdd 17_3/a_26_538# 3.79359f
C30 GND 17_28/a_62_902# 2.79216f
C31 GND 17_3/DI 4.11066f
C32 GND 17_9/DIB 6.35733f
C33 GND 17_13/OEN 4.46481f
C34 Vdd 17_13/DO 3.11769f
C35 17_4/a_420_786# p_b 2.95776f
C36 GND 17_11/DIB 6.35733f
C37 Vdd 17_28/DIB 6.39135f
C38 GND 17_28/a_58_538# 3.79746f
C39 17_7/a_62_902# p_h 6.99264f
C40 GND 17_19/a_62_902# 2.79216f
C41 p_b 17_4/a_62_82# 8.056081f
C42 17_14/w_40_1480# 17_14/DATA 66.6688f
C43 Vdd 17_2/a_26_538# 3.76551f
C44 GND p_a 0.100362p
C45 Vdd 17_19/DIB 6.39135f
C46 GND 17_19/a_58_538# 3.79746f
C47 GND 17_17/a_62_902# 2.79216f
C48 Vdd 17_15/a_26_538# 3.76551f
C49 GND 17_15/DATA 0.100362p
C50 Vdd 17_29/a_58_538# 6.72912f
C51 GND 17_8/DIB 6.35733f
C52 GND 17_12/OEN 4.46481f
C53 Vdd 17_12/DO 3.11769f
C54 Vdd 17_17/DIB 6.39135f
C55 GND 17_17/a_58_538# 3.79746f
C56 GND 17_15/DI 4.11066f
C57 17_3/w_40_1480# p_i 66.6688f
C58 17_14/a_420_786# 17_14/DATA 2.95776f
C59 GND 17_31/OEN 4.46481f
C60 Vdd 17_31/DO 3.11769f
C61 17_20/a_252_786# 17_20/DATA 3.00456f
C62 Vdd 17_0/a_26_538# 3.76551f
C63 GND 17_0/DATA 0.100362p
C64 GND 17_0/DI 4.11066f
C65 GND 17_27/a_62_902# 2.79216f
C66 Vdd 17_25/a_26_538# 3.76551f
C67 GND 17_25/DATA 0.100362p
C68 17_32/w_40_1480# 17_32/DATA 66.6688f
C69 GND 17_7/DIB 6.35733f
C70 17_3/a_420_786# p_i 2.95776f
C71 Vdd 17_27/DIB 6.39135f
C72 GND 17_27/a_58_538# 3.79746f
C73 Vdd 17_35/a_26_538# 3.76551f
C74 GND 17_35/DATA 0.100362p
C75 17_6/a_62_902# p_c 6.99264f
C76 GND 17_25/DI 4.11066f
C77 p_i 17_3/a_62_82# 8.056081f
C78 GND 17_35/DI 4.11066f
C79 GND 17_20/OEN 4.46481f
C80 Vdd 17_20/DO 3.11769f
C81 Vdd 17_1/a_26_538# 3.76551f
C82 GND 17_1/DATA 0.100362p
C83 GND 17_29/DO 4.38615f
C84 17_32/a_420_786# 17_32/DATA 2.95776f
C85 GND 17_16/a_62_902# 2.79216f
C86 GND 17_1/DI 4.11066f
C87 GND 17_6/DIB 6.35733f
C88 Vdd 17_32/DATA 0.111498p
C89 17_32/DATA 17_32/a_62_82# 8.056081f
C90 Vdd 17_16/DIB 6.39135f
C91 GND 17_16/a_58_538# 3.79746f
C92 Vdd 17_34/a_26_538# 3.76551f
C93 GND 17_34/DATA 0.100362p
C94 Vdd GND 5.46408p
C95 17_2/w_40_1480# p_a 66.6688f
C96 Vdd 17_32/DI 3.31488f
C97 GND 17_32/a_62_82# 48.660957f
C98 GND b 4.32666f
C99 Vdd a 4.34502f
C100 GND 17_34/DI 4.11066f
C101 GND 17_30/OEN 4.46481f
C102 Vdd 17_30/DO 3.11769f
C103 17_30/a_252_786# 17_30/DATA 3.00456f
C104 GND 17_26/a_62_902# 2.79216f
C105 17_15/w_40_1480# 17_15/DATA 66.6688f
C106 Vdd 17_33/a_62_902# 51.916096f
C107 17_21/w_40_1480# 17_21/DATA 66.6688f
C108 GND 17_5/DIB 6.35733f
C109 Vdd 17_21/DATA 0.111498p
C110 17_2/a_420_786# p_a 2.95776f
C111 Vdd 17_26/DIB 6.39135f
C112 GND 17_26/a_58_538# 3.79746f
C113 Vdd 17_24/a_26_538# 3.76551f
C114 GND 17_24/DATA 0.100362p
C115 17_5/a_62_902# p_d 6.99264f
C116 GND 17_33/DO 4.38615f
C117 Vdd 17_33/a_58_538# 6.72912f
C118 Vdd 17_21/DI 3.31488f
C119 GND 17_21/a_62_82# 48.660957f
C120 p_a 17_2/a_62_82# 8.056081f
C121 Vdd c 4.95882f
C122 GND 17_24/DI 4.11066f
C123 17_15/a_420_786# 17_15/DATA 2.95776f
C124 17_21/a_420_786# 17_21/DATA 2.95776f
C125 Vdd 17_22/a_62_902# 51.916096f
C126 Vdd 17_10/DATA 0.111498p
C127 GND 17_4/DIB 6.35733f
C128 17_15/DATA 17_15/a_62_82# 8.056081f
C129 17_29/DATA 17_29/a_420_786# 2.95776f
C130 17_21/DATA 17_21/a_62_82# 8.056081f
C131 Vdd 17_23/a_26_538# 3.76551f
C132 GND 17_23/DATA 0.100362p
C133 GND 17_22/DO 4.38615f
C134 Vdd 17_22/a_58_538# 6.72912f
C135 17_0/w_40_1480# 17_0/DATA 66.6688f
C136 GND 17_18/OEN 4.46481f
C137 Vdd 17_18/DO 3.11769f
C138 Vdd 17_10/DI 3.31488f
C139 GND 17_10/a_62_82# 48.660957f
C140 17_14/m3_n72_n22# GND 32.52166f
C141 GND 17_23/DI 4.11066f
C142 Vdd 17_9/a_62_902# 51.916096f
C143 17_25/w_40_1480# 17_25/DATA 66.6688f
C144 Vdd 17_11/a_62_902# 51.916096f
C145 17_10/w_40_1480# 17_10/DATA 66.6688f
C146 GND 17_3/DIB 6.35733f
C147 GND 17_9/DO 4.38615f
C148 Vdd 17_9/a_58_538# 6.72912f
C149 17_0/a_420_786# 17_0/DATA 2.95776f
C150 Vdd 17_13/a_26_538# 3.76551f
C151 GND 17_13/DATA 0.100362p
C152 17_4/a_62_902# p_b 6.99264f
C153 GND 17_28/OEN 4.46481f
C154 Vdd 17_28/DO 3.11769f
C155 GND 17_11/DO 4.38615f
C156 Vdd 17_11/a_58_538# 6.72912f
C157 17_0/DATA 17_0/a_62_82# 8.056081f
C158 17_35/w_40_1480# 17_35/DATA 66.6688f
C159 GND 17_13/DI 4.11066f
C160 17_25/a_420_786# 17_25/DATA 2.95776f
C161 Vdd 17_8/a_62_902# 51.916096f
C162 GND 17_19/OEN 4.46481f
C163 Vdd 17_19/DO 3.11769f
C164 17_10/a_420_786# 17_10/DATA 2.95776f
C165 GND 17_2/DIB 6.35733f
C166 17_18/a_252_786# 17_18/DATA 3.00456f
C167 17_25/DATA 17_25/a_62_82# 8.056081f
C168 GND 17_8/DO 4.38615f
C169 Vdd 17_8/a_58_538# 6.72912f
C170 17_10/DATA 17_10/a_62_82# 8.056081f
C171 Vdd 17_12/a_26_538# 3.76551f
C172 GND 17_12/DATA 0.100362p
C173 GND 17_17/OEN 4.46481f
C174 Vdd 17_17/DO 3.11769f
C175 17_35/a_420_786# 17_35/DATA 2.95776f
C176 17_1/w_40_1480# 17_1/DATA 66.6688f
C177 GND 17_15/DIB 6.35733f
C178 17_14/a_62_902# 17_14/DATA 6.99264f
C179 GND 17_12/DI 4.11066f
C180 17_35/DATA 17_35/a_62_82# 8.056081f
C181 Vdd 17_31/a_26_538# 3.76551f
C182 GND 17_31/DATA 0.100362p
C183 Vdd 17_29/a_26_538# 3.76551f
C184 Vdd 17_7/a_62_902# 51.916096f
C185 GND 17_31/DI 4.11066f
C186 GND 17_0/DIB 6.35733f
C187 Vdd 17_7/a_58_538# 6.72912f
C188 17_1/a_420_786# 17_1/DATA 2.95776f
C189 17_3/a_62_902# p_i 6.99264f
C190 GND 17_27/OEN 4.46481f
C191 Vdd 17_27/DO 3.11769f
C192 17_29/DATA 17_29/a_62_82# 8.056081f
C193 GND 17_25/DIB 6.35733f
C194 17_34/w_40_1480# 17_34/DATA 66.6688f
C195 17_1/DATA 17_1/a_62_82# 8.056081f
C196 GND 17_35/DIB 6.35733f
C197 Vdd 17_20/a_26_538# 3.76551f
C198 GND 17_20/DATA 0.100362p
C199 Vdd 17_6/a_62_902# 51.916096f
C200 GND 17_20/DI 4.11066f
C201 17_32/a_62_902# 17_32/DATA 6.99264f
C202 GND 17_1/DIB 6.35733f
C203 17_28/a_252_786# 17_28/DATA 3.00456f
C204 GND 17_32/a_62_902# 2.79216f
C205 GND 17_6/DO 4.38615f
C206 Vdd 17_6/a_58_538# 6.72912f
C207 GND 17_16/OEN 4.46481f
C208 Vdd 17_16/DO 3.11769f
C209 GND 17_29/a_62_902# 2.79216f
C210 17_34/a_420_786# 17_34/DATA 2.95776f
C211 Vdd 17_32/DIB 6.39135f
C212 GND 17_32/a_58_538# 3.79746f
C213 Vdd 17_29/DI 3.31488f
C214 GND 19_1/w_40_1480# 66.6688f
C215 GND 17_34/DIB 6.35733f
C216 17_34/DATA 17_34/a_62_82# 8.056081f
C217 Vdd 17_30/a_26_538# 3.76551f
C218 GND 17_30/DATA 0.100362p
C219 Vdd 17_5/a_62_902# 51.916096f
C220 GND 17_30/DI 4.11066f
C221 17_19/a_252_786# 17_19/DATA 3.00456f
C222 GND 17_5/DO 4.38615f
C223 Vdd 17_5/a_58_538# 6.72912f
C224 GND 17_21/a_62_902# 2.79216f
C225 17_2/a_62_902# p_a 6.99264f
C226 GND 17_26/OEN 4.46481f
C227 Vdd 17_26/DO 3.11769f
C228 GND 17_33/a_26_538# 3.75903f
C229 Vdd 17_21/DIB 6.39135f
C230 GND 17_21/a_58_538# 3.79746f
C231 17_24/w_40_1480# 17_24/DATA 66.6688f
C232 Vdd 17_29/DIB 6.39135f
C233 GND 17_24/DIB 6.35733f
C234 GND 17_33/m3_n72_n22# 32.52166f
C235 Vdd 17_4/a_62_902# 51.916096f
C236 17_15/a_62_902# 17_15/DATA 6.99264f
C237 17_21/a_62_902# 17_21/DATA 6.99264f
C238 17_17/a_252_786# 17_17/DATA 3.00456f
C239 GND 17_4/DO 4.38615f
C240 Vdd 17_4/a_58_538# 6.72912f
C241 17_33/a_252_786# 17_33/DATA 3.00456f
C242 GND 17_10/a_62_902# 2.79216f
C243 17_24/a_420_786# 17_24/DATA 2.95776f
C244 GND 17_22/a_26_538# 3.75903f
C245 Vdd 17_18/a_26_538# 3.76551f
C246 GND 17_18/DATA 0.100362p
C247 Vdd 17_10/DIB 6.39135f
C248 GND 17_10/a_58_538# 3.79746f
C249 17_14/DI Vdd 3.31488f
C250 17_14/a_62_82# GND 48.660957f
C251 17_14/a_62_902# Vdd 51.916096f
C252 17_24/DATA 17_24/a_62_82# 8.056081f
C253 GND 17_23/DIB 6.35733f
C254 GND 17_22/m3_n72_n22# 32.52166f
C255 GND 17_18/DI 4.11066f
C256 17_14/DO GND 4.38615f
C257 Vdd 17_3/a_62_902# 51.916096f
C258 Vdd 18_1/w_40_1480# 66.6688f
C259 Vdd 17_3/a_58_538# 6.72912f
C260 GND 17_9/a_26_538# 3.75903f
C261 17_0/a_62_902# 17_0/DATA 6.99264f
C262 GND 17_11/a_26_538# 3.75903f
C263 Vdd 17_28/a_26_538# 3.76551f
C264 GND 17_28/DATA 0.100362p
C265 17_23/w_40_1480# 17_23/DATA 66.6688f
C266 GND 17_9/m3_n72_n22# 32.52166f
C267 Vdd 17_29/DATA 0.111498p
C268 GND 17_13/DIB 6.35733f
C269 GND 17_28/DI 4.11066f
C270 GND 17_11/m3_n72_n22# 32.52166f
C271 Vdd 17_2/a_62_902# 51.916096f
C272 17_25/a_62_902# 17_25/DATA 6.99264f
C273 Vdd 17_19/a_26_538# 3.76551f
C274 GND 17_19/DATA 0.100362p
C275 17_10/a_62_902# 17_10/DATA 6.99264f
C276 17_27/a_252_786# 17_27/DATA 3.00456f
C277 GND 17_2/DO 4.38615f
C278 Vdd 17_2/a_58_538# 6.72912f
C279 17_22/a_252_786# 17_22/DATA 3.00456f
C280 Vdd 17_15/a_62_902# 51.916096f
C281 GND 17_8/a_26_538# 3.75903f
C282 GND 17_19/DI 4.11066f
C283 17_23/a_420_786# 17_23/DATA 2.95776f
C284 17_14/a_58_538# Vdd 6.72912f
C285 Vdd 17_17/a_26_538# 3.76551f
C286 GND 17_17/DATA 0.100362p
C287 17_35/a_62_902# 17_35/DATA 6.99264f
C288 GND 17_15/DO 4.38615f
C289 Vdd 17_15/a_58_538# 6.72912f
C290 GND 17_8/m3_n72_n22# 32.52166f
C291 17_23/DATA 17_23/a_62_82# 8.056081f
C292 GND 17_12/DIB 6.35733f
C293 GND 17_17/DI 4.11066f
C294 Vdd 17_0/a_62_902# 51.916096f
C295 GND 17_31/DIB 6.35733f
C296 GND 17_0/DO 4.38615f
C297 Vdd 17_0/a_58_538# 6.72912f
C298 Vdd 17_25/a_62_902# 51.916096f
C299 GND 17_7/a_26_538# 3.75903f
C300 17_1/a_62_902# 17_1/DATA 6.99264f
C301 Vdd 17_27/a_26_538# 3.76551f
C302 GND 17_27/DATA 0.100362p
C303 Vdd 17_35/a_62_902# 51.916096f
C304 GND 17_25/DO 4.38615f
C305 Vdd 17_25/a_58_538# 6.72912f
C306 17_13/w_40_1480# 17_13/DATA 66.6688f
C307 GND 17_7/m3_n72_n22# 32.52166f
C308 GND 17_27/DI 4.11066f
C309 GND 17_35/DO 4.38615f
C310 Vdd 17_35/a_58_538# 6.72912f
C311 17_9/a_252_786# 17_9/DATA 3.00456f
C312 Vdd 17_1/a_62_902# 51.916096f
C313 GND 17_20/DIB 6.35733f
C314 17_16/a_252_786# 17_16/DATA 3.00456f
C315 GND 17_1/DO 4.38615f
C316 Vdd 17_1/a_58_538# 6.72912f
C317 17_11/a_252_786# 17_11/DATA 3.00456f
C318 GND 17_6/a_26_538# 3.78711f
C319 17_13/a_420_786# 17_13/DATA 2.95776f
C320 Vdd 17_16/a_26_538# 3.76551f
C321 GND 17_16/DATA 0.100362p
C322 17_34/a_62_902# 17_34/DATA 6.99264f
C323 Vdd 17_34/a_62_902# 51.916096f
C324 GND 17_32/OEN 4.46481f
C325 Vdd 17_32/DO 3.11769f
C326 GND 17_6/m3_n72_n22# 33.6463f
C327 17_13/DATA 17_13/a_62_82# 8.056081f
C328 GND 17_16/DI 4.11066f
C329 GND 17_34/DO 4.38615f
C330 Vdd 17_34/a_58_538# 6.72912f
C331 GND i 4.76415f
C332 GND 17_30/DIB 6.35733f
C333 GND 17_5/a_26_538# 3.78711f
C334 Vdd 17_26/a_26_538# 3.76551f
C335 GND 17_26/DATA 0.100362p
C336 Vdd 17_24/a_62_902# 51.916096f
C337 17_12/w_40_1480# 17_12/DATA 66.6688f
C338 Vdd 17_33/DATA 0.111498p
C339 GND 17_5/m3_n72_n22# 33.2755f
C340 GND 17_21/OEN 4.46481f
C341 Vdd 17_21/DO 3.11769f
C342 GND 17_26/DI 4.11066f
C343 GND 17_24/DO 4.38615f
C344 Vdd 17_24/a_58_538# 6.72912f
C345 Vdd 17_33/DI 3.31488f
C346 GND 17_33/a_62_82# 48.660957f
C347 17_8/a_252_786# 17_8/DATA 3.00456f
C348 GND h 4.65615f
C349 17_26/a_252_786# 17_26/DATA 3.00456f
C350 GND 17_4/a_26_538# 3.78711f
C351 17_31/w_40_1480# 17_31/DATA 66.6688f
C352 17_12/a_420_786# 17_12/DATA 2.95776f
C353 17_24/a_62_902# 17_24/DATA 6.99264f
C354 Vdd 17_23/a_62_902# 51.916096f
C355 Vdd 17_22/DATA 0.111498p
C356 GND 17_4/m3_n72_n22# 33.2755f
C357 GND 17_10/OEN 4.46481f
C358 Vdd 17_10/DO 3.11769f
C359 17_14/DIB Vdd 6.39135f
C360 17_12/DATA 17_12/a_62_82# 8.056081f
C361 GND d 5.21766f
C362 GND 17_23/DO 4.38615f
C363 Vdd 17_23/a_58_538# 6.72912f
C364 Vdd 17_22/DI 3.31488f
C365 GND 17_22/a_62_82# 48.660957f
C366 GND 17_18/DIB 6.35733f
C367 17_14/a_26_538# GND 3.75903f
C368 17_31/a_420_786# 17_31/DATA 2.95776f
C369 GND 17_3/a_26_538# 3.75903f
C370 Vdd 17_9/DATA 0.111498p
C371 17_31/DATA 17_31/a_62_82# 8.056081f
C372 Vdd 17_13/a_62_902# 51.916096f
C373 Vdd 17_11/DATA 0.111498p
C374 GND 17_3/m3_n72_n22# 32.52166f
C375 Vdd 17_9/DI 3.31488f
C376 GND 17_9/a_62_82# 48.660957f
C377 17_29/DATA 17_29/a_62_902# 6.99264f
C378 GND 17_13/DO 4.38615f
C379 Vdd 17_13/a_58_538# 6.72912f
C380 Vdd 17_11/DI 3.31488f
C381 GND 17_11/a_62_82# 48.660957f
C382 GND 17_28/DIB 6.35733f
C383 17_7/a_252_786# p_h 3.00456f
C384 GND 17_2/a_26_538# 3.78711f
C385 17_20/w_40_1480# 17_20/DATA 66.6688f
C386 GND 17_19/DIB 6.35733f
C387 Vdd 17_8/DATA 0.111498p
C388 17_23/a_62_902# 17_23/DATA 6.99264f
C389 Vdd 17_12/a_62_902# 51.916096f
C390 GND 17_2/m3_n72_n22# 33.2755f
C391 GND 17_15/a_26_538# 3.75903f
C392 GND 17_29/a_58_538# 3.79746f
C393 Vdd 17_8/DI 3.31488f
C394 GND 17_8/a_62_82# 48.660957f
C395 GND 17_12/DO 4.38615f
C396 Vdd 17_12/a_58_538# 6.72912f
C397 GND 17_17/DIB 6.35733f
C398 Vdd 17_31/a_62_902# 51.916096f
C399 GND 17_15/m3_n72_n22# 32.52166f
C400 GND 17_31/DO 4.38615f
C401 Vdd 17_31/a_58_538# 6.72912f
C402 17_20/a_420_786# 17_20/DATA 2.95776f
C403 GND 17_0/a_26_538# 3.78711f
C404 Vdd p_h 0.111498p
C405 17_20/DATA 17_20/a_62_82# 8.056081f
C406 GND 17_0/m3_n72_n22# 34.6831f
C407 GND 17_25/a_26_538# 3.75903f
C408 Vdd 17_7/DI 3.31488f
C409 GND 17_7/a_62_82# 48.660957f
C410 GND 17_27/DIB 6.35733f
C411 GND 17_35/a_26_538# 3.75903f
C412 17_6/a_252_786# p_c 3.00456f
C413 GND 17_26/m3_n72_n22# 61.8451f
C414 Vdd 17_20/a_62_902# 51.916096f
C415 GND 17_35/m3_n72_n22# 32.52166f
C416 GND 17_20/DO 4.38615f
C417 Vdd 17_20/a_58_538# 6.72912f
C418 GND 17_1/a_26_538# 3.75903f
C419 17_30/w_40_1480# 17_30/DATA 66.6688f
C420 Vdd p_c 0.111498p
C421 GND 17_29/m3_n72_n22# 32.52166f
C422 17_13/a_62_902# 17_13/DATA 6.99264f
C423 GND 17_1/m3_n72_n22# 32.52166f
C424 GND 17_6/a_62_82# 48.660957f
C425 Vdd 17_32/a_26_538# 3.76551f
C426 GND 17_32/DATA 0.100362p
C427 GND 17_16/DIB 6.35733f
C428 GND 17_34/a_26_538# 3.75903f
C429 Vdd 17_30/a_62_902# 51.916096f
C430 GND a 4.32666f
C431 GND 17_32/DI 4.11066f
C432 GND 17_34/m3_n72_n22# 33.929264f
C433 GND 17_30/DO 4.38615f
C434 Vdd 17_30/a_58_538# 6.72912f
C435 17_30/a_420_786# 17_30/DATA 2.95776f
C436 Vdd p_d 0.111498p
C437 17_30/DATA 17_30/a_62_82# 8.056081f
C438 GND 17_33/a_62_902# 2.79216f
C439 GND 17_5/a_62_82# 48.660957f
C440 Vdd 17_21/a_26_538# 3.76551f
C441 GND 17_21/DATA 0.100362p
C442 GND 17_26/DIB 6.35733f
C443 GND 17_24/a_26_538# 3.75903f
C444 17_5/a_252_786# p_d 3.00456f
C445 Vdd 17_33/DIB 6.39135f
C446 GND 17_33/a_58_538# 3.79746f
C447 GND 17_21/DI 4.11066f
C448 GND c 4.32666f
C449 GND 17_24/m3_n72_n22# 32.52166f
C450 Vdd p_b 0.111498p
C451 17_12/a_62_902# 17_12/DATA 6.99264f
C452 GND 17_22/a_62_902# 2.79216f
C453 GND 17_4/a_62_82# 48.660957f
C454 Vdd 17_18/a_62_902# 51.916096f
C455 Vdd 17_10/a_26_538# 3.76551f
C456 GND 17_10/DATA 0.100362p
C457 GND 17_23/a_26_538# 3.75903f
C458 GND 17_18/DO 4.38615f
C459 Vdd 17_18/a_58_538# 6.72912f
C460 Vdd 17_22/DIB 6.39135f
C461 GND 17_22/a_58_538# 3.79746f
C462 GND 17_10/DI 4.11066f
C463 17_14/DATA Vdd 0.111498p
C464 GND 17_23/m3_n72_n22# 32.52166f
C465 17_29/DATA 17_29/w_40_1480# 66.6688f
C466 17_31/a_62_902# 17_31/DATA 6.99264f
C467 Vdd p_i 0.111498p
C468 GND 17_9/a_62_902# 2.79216f
C469 Vdd 17_28/a_62_902# 51.916096f
C470 GND 17_11/a_62_902# 2.79216f
C471 Vdd 17_3/DI 3.31488f
C472 GND 17_3/a_62_82# 48.660957f
C473 Vdd 17_9/DIB 6.39135f
C474 GND 17_9/a_58_538# 3.79746f
C475 17_18/w_40_1480# 17_18/DATA 66.6688f
C476 GND 17_13/a_26_538# 3.75903f
C477 17_4/a_252_786# p_b 3.00456f
C478 Vdd 17_11/DIB 6.39135f
C479 GND 17_11/a_58_538# 3.79746f
C480 GND 17_28/DO 4.38615f
C481 Vdd 17_28/a_58_538# 6.72912f
C482 GND 17_13/m3_n72_n22# 32.78878f
C483 Vdd 17_19/a_62_902# 51.916096f
C484 Vdd p_a 0.111498p
C485 GND 17_19/DO 4.38615f
C486 Vdd 17_19/a_58_538# 6.72912f
C487 GND 17_8/a_62_902# 2.79216f
C488 Vdd 17_17/a_62_902# 51.916096f
C489 GND 17_2/a_62_82# 48.660957f
C490 17_18/a_420_786# 17_18/DATA 2.95776f
C491 Vdd 17_15/DATA 0.111498p
C492 Vdd 17_8/DIB 6.39135f
C493 GND 17_8/a_58_538# 3.79746f
C494 GND 17_12/a_26_538# 3.75903f
C495 GND 17_17/DO 4.38615f
C496 Vdd 17_17/a_58_538# 6.72912f
C497 17_18/DATA 17_18/a_62_82# 8.056081f
C498 Vdd 17_15/DI 3.31488f
C499 GND 17_15/a_62_82# 48.660957f
C500 17_14/a_252_786# 17_14/DATA 3.00456f
C501 GND 17_12/m3_n72_n22# 32.78878f
C502 GND 17_31/a_26_538# 3.75903f
C503 GND 17_29/a_26_538# 3.75903f
C504 17_20/a_62_902# 17_20/DATA 6.99264f
C505 Vdd 17_0/DATA 0.111498p
C506 GND 17_7/a_62_902# 2.79216f
C507 GND 17_31/m3_n72_n22# 32.52166f
C508 Vdd 17_27/a_62_902# 51.916096f
C509 Vdd 17_0/DI 3.31488f
C510 GND 17_0/a_62_82# 48.660957f
C511 Vdd 17_25/DATA 0.111498p
C512 Vdd 17_7/DIB 6.39135f
C513 GND 17_7/a_58_538# 3.79746f
C514 17_28/w_40_1480# 17_28/DATA 66.6688f
C515 17_3/a_252_786# p_i 3.00456f
C516 GND 17_27/DO 4.38615f
C517 Vdd 17_27/a_58_538# 6.72912f
C518 Vdd 17_35/DATA 0.111498p
C519 Vdd 17_25/DI 3.31488f
C520 GND 17_25/a_62_82# 48.660957f
C521 Vdd 17_35/DI 3.31488f
C522 GND 17_35/a_62_82# 48.660957f
C523 GND 17_20/a_26_538# 3.75903f
C524 Vdd 17_1/DATA 0.111498p
C525 GND 17_6/a_62_902# 2.79216f
C526 Vdd 17_29/DO 3.11769f
C527 GND 17_20/m3_n72_n22# 32.52166f
C528 17_32/a_252_786# 17_32/DATA 3.00456f
C529 Vdd 17_1/DI 3.31488f
C530 GND 17_1/a_62_82# 48.660957f
C531 17_28/a_420_786# 17_28/DATA 2.95776f
C532 Vdd 17_16/a_62_902# 51.916096f
C533 Vdd 17_6/DIB 6.39135f
C534 GND 17_6/a_58_538# 3.79746f
C535 GND 17_16/DO 4.38615f
C536 Vdd 17_16/a_58_538# 6.72912f
C537 Vdd 17_34/DATA 0.111498p
C538 17_28/DATA 17_28/a_62_82# 8.056081f
C539 GND 17_32/DIB 6.35733f
C540 GND 17_29/DI 4.11066f
C541 Vdd b 3.6576f
C542 Vdd 17_34/DI 3.31488f
C543 GND 17_34/a_62_82# 48.660957f
C544 17_30/a_62_902# 17_30/DATA 6.99264f
C545 GND 17_30/a_26_538# 3.75903f
C546 GND 17_5/a_62_902# 2.79216f
C547 GND 17_30/m3_n72_n22# 32.89246f
C548 Vdd 17_26/a_62_902# 51.916096f
C549 17_19/a_420_786# 17_19/DATA 2.95776f
C550 Vdd 17_5/DIB 6.39135f
C551 GND 17_5/a_58_538# 3.79746f
C552 17_17/w_40_1480# 17_17/DATA 66.6688f
C553 17_2/a_252_786# p_a 3.00456f
C554 17_33/w_40_1480# 17_33/DATA 66.6688f
C555 GND 17_26/DO 4.38615f
C556 Vdd 17_26/a_58_538# 6.72912f
C557 Vdd 17_24/DATA 0.111498p
C558 GND 17_33/OEN 4.46481f
C559 Vdd 17_33/DO 3.11769f
C560 17_19/DATA 17_19/a_62_82# 8.056081f
C561 GND 17_21/DIB 6.35733f
C562 GND 17_29/DIB 6.35733f
C563 Vdd 17_24/DI 3.31488f
C564 GND 17_24/a_62_82# 48.660957f
C565 GND 17_29/OEN 4.46481f
C566 GND 17_4/a_62_902# 2.79216f
C567 17_15/a_252_786# 17_15/DATA 3.00456f
C568 17_21/a_252_786# 17_21/DATA 3.00456f
C569 17_17/a_420_786# 17_17/DATA 2.95776f
C570 Vdd 17_4/DIB 6.39135f
C571 GND 17_4/a_58_538# 3.79746f
C572 17_33/a_420_786# 17_33/DATA 2.95776f
C573 Vdd 17_23/DATA 0.111498p
C574 17_17/DATA 17_17/a_62_82# 8.056081f
C575 GND 17_22/OEN 4.46481f
C576 Vdd 17_22/DO 3.11769f
C577 GND 17_18/a_26_538# 3.75903f
C578 17_33/DATA 17_33/a_62_82# 8.056081f
C579 GND 17_10/DIB 6.35733f
C580 17_14/a_62_902# GND 2.79216f
C581 17_14/DI GND 4.11066f
C582 Vdd 17_23/DI 3.31488f
C583 GND 17_23/a_62_82# 48.660957f
C584 GND 17_18/m3_n72_n22# 32.52166f
C585 GND 17_3/a_62_902# 2.79216f
C586 17_29/DATA 17_29/a_252_786# 3.00456f
C587 Vdd 17_3/DIB 6.39135f
C588 GND 17_3/a_58_538# 3.79746f
C589 17_27/w_40_1480# 17_27/DATA 66.6688f
C590 GND 17_9/OEN 4.46481f
C591 Vdd 17_9/DO 3.11769f
C592 17_0/a_252_786# 17_0/DATA 3.00456f
C593 17_22/w_40_1480# 17_22/DATA 66.6688f
C594 Vdd 17_13/DATA 0.111498p
C595 GND 17_28/a_26_538# 3.75903f
C596 GND 17_11/OEN 4.46481f
C597 Vdd 17_11/DO 3.11769f
C598 GND 17_29/DATA 0.100362p
C599 Vdd 17_13/DI 3.31488f
C600 GND 17_13/a_62_82# 48.660957f
C601 GND 17_28/m3_n72_n22# 32.52166f
C602 GND 17_2/a_62_902# 2.79216f
C603 17_25/a_252_786# 17_25/DATA 3.00456f
C604 GND 17_19/a_26_538# 3.75903f
C605 17_10/a_252_786# 17_10/DATA 3.00456f
C606 17_27/a_420_786# 17_27/DATA 2.95776f
C607 Vdd 17_2/DIB 6.39135f
C608 GND 17_2/a_58_538# 3.79746f
C609 17_18/a_62_902# 17_18/DATA 6.99264f
C610 17_22/a_420_786# 17_22/DATA 2.95776f
C611 GND 17_19/m3_n72_n22# 32.52166f
C612 GND 17_15/a_62_902# 2.79216f
C613 GND 17_8/OEN 4.46481f
C614 Vdd 17_8/DO 3.11769f
C615 Vdd 17_12/DATA 0.111498p
C616 17_27/DATA 17_27/a_62_82# 8.056081f
C617 17_14/a_58_538# GND 3.79746f
C618 GND 17_17/a_26_538# 3.75903f
C619 17_35/a_252_786# 17_35/DATA 3.00456f
C620 Vdd 17_15/DIB 6.39135f
C621 GND 17_15/a_58_538# 3.79746f
C622 17_22/DATA 17_22/a_62_82# 8.056081f
C623 17_14/DATA 17_14/a_62_82# 8.056081f
C624 Vdd 17_12/DI 3.31488f
C625 GND 17_12/a_62_82# 48.660957f
C626 GND 17_17/m3_n72_n22# 32.52166f
C627 Vdd 17_31/DATA 0.111498p
C628 GND 17_0/a_62_902# 2.79216f
C629 17_9/w_40_1480# 17_9/DATA 66.6688f
C630 Vdd 17_31/DI 3.31488f
C631 GND 17_31/a_62_82# 48.660957f
C632 Vdd 17_0/DIB 6.39135f
C633 GND 17_0/a_58_538# 3.79746f
C634 GND 17_25/a_62_902# 2.79216f
C635 17_16/w_40_1480# 17_16/DATA 66.6688f
C636 17_1/a_252_786# 17_1/DATA 3.00456f
C637 17_11/w_40_1480# 17_11/DATA 66.6688f
C638 GND 17_27/a_26_538# 3.75903f
C639 GND 17_35/a_62_902# 2.79216f
C640 Vdd 17_25/DIB 6.39135f
C641 GND 17_25/a_58_538# 3.79746f
C642 17_19/w_40_1480# 17_19/DATA 66.6688f
C643 GND 17_27/m3_n72_n22# 32.52166f
C644 Vdd 17_35/DIB 6.39135f
C645 GND 17_35/a_58_538# 3.79746f
C646 Vdd 17_20/DATA 0.111498p
C647 17_9/a_420_786# 17_9/DATA 2.95776f
C648 GND 17_1/a_62_902# 2.79216f
C649 Vdd 17_20/DI 3.31488f
C650 GND 17_20/a_62_82# 48.660957f
C651 17_16/a_420_786# 17_16/DATA 2.95776f
C652 17_9/DATA 17_9/a_62_82# 8.056081f
C653 17_11/a_420_786# 17_11/DATA 2.95776f
C654 Vdd 17_1/DIB 6.39135f
C655 GND 17_1/a_58_538# 3.79746f
C656 17_28/a_62_902# 17_28/DATA 6.99264f
C657 Vdd 17_6/DO 3.11769f
C658 Vdd 17_32/a_62_902# 51.916096f
C659 17_16/DATA 17_16/a_62_82# 8.056081f
C660 Vdd 17_29/a_62_902# 51.916096f
C661 GND 17_16/a_26_538# 3.75903f
C662 GND 17_34/a_62_902# 2.79216f
C663 17_34/a_252_786# 17_34/DATA 3.00456f
C664 17_11/DATA 17_11/a_62_82# 8.056081f
C665 GND 17_32/DO 4.38615f
C666 Vdd 17_32/a_58_538# 6.72912f
C667 GND 17_16/m3_n72_n22# 32.52166f
C668 Vdd 17_34/DIB 6.39135f
C669 GND 17_34/a_58_538# 3.79746f
C670 Vdd 17_30/DATA 0.111498p
C671 17_8/w_40_1480# 17_8/DATA 66.6688f
C672 Vdd 17_30/DI 3.31488f
C673 GND 17_30/a_62_82# 48.660957f
C674 17_19/a_62_902# 17_19/DATA 6.99264f
C675 Vdd 17_5/DO 3.11769f
C676 17_26/w_40_1480# 17_26/DATA 66.6688f
C677 Vdd 17_21/a_62_902# 51.916096f
C678 GND 17_26/a_26_538# 3.75903f
C679 GND 17_24/a_62_902# 2.79216f
C680 Vdd 17_33/a_26_538# 3.76551f
C681 GND 17_33/DATA 0.100362p
C682 GND 17_21/DO 4.38615f
C683 Vdd 17_21/a_58_538# 6.72912f
C684 Vdd 17_24/DIB 6.39135f
C685 GND 17_24/a_58_538# 3.79746f
C686 GND 17_33/DI 4.11066f
C687 17_8/a_420_786# 17_8/DATA 2.95776f
C688 17_26/a_420_786# 17_26/DATA 2.95776f
C689 17_8/DATA 17_8/a_62_82# 8.056081f
C690 GND 19_0/w_40_1480# 66.6688f
C691 17_17/a_62_902# 17_17/DATA 6.99264f
C692 Vdd 17_4/DO 3.11769f
C693 17_33/a_62_902# 17_33/DATA 6.99264f
C694 Vdd 17_10/a_62_902# 51.916096f
C695 17_26/DATA 17_26/a_62_82# 8.056081f
C696 17_24/a_252_786# 17_24/DATA 3.00456f
C697 GND 17_23/a_62_902# 2.79216f
C698 Vdd 17_22/a_26_538# 3.76551f
C699 GND 17_22/DATA 0.100362p
C700 Vdd 17_18/DATA 0.111498p
C701 GND 17_10/DO 4.38615f
C702 Vdd 17_10/a_58_538# 6.72912f
C703 17_14/DIB GND 6.35733f
C704 Vdd 17_23/DIB 6.39135f
C705 GND 17_23/a_58_538# 3.79746f
C706 GND 17_22/DI 4.11066f
C707 Vdd 17_18/DI 3.31488f
C708 GND 17_18/a_62_82# 48.660957f
C709 17_14/OEN GND 4.46481f
C710 17_14/DO Vdd 3.11769f
C711 17_7/w_40_1480# p_h 66.6688f
C712 Vdd 17_9/a_26_538# 3.76551f
C713 GND 17_9/DATA 0.100362p
C714 GND 17_13/a_62_902# 2.79216f
C715 Vdd 17_11/a_26_538# 3.76551f
C716 GND 17_11/DATA 0.100362p
C717 Vdd 17_28/DATA 0.111498p
C718 GND 17_9/DI 4.11066f
C719 Vdd 17_13/DIB 6.39135f
C720 GND 17_13/a_58_538# 3.79746f
C721 GND 17_11/DI 4.11066f
C722 Vdd 17_28/DI 3.31488f
C723 GND 17_28/a_62_82# 48.660957f
C724 17_7/a_420_786# p_h 2.95776f
C725 Vdd 17_19/DATA 0.111498p
C726 p_h 17_7/a_62_82# 8.056081f
C727 17_27/a_62_902# 17_27/DATA 6.99264f
C728 17_22/a_62_902# 17_22/DATA 6.99264f
C729 Vdd 17_2/DO 3.11769f
C730 Vdd 17_19/DI 3.31488f
C731 GND 17_19/a_62_82# 48.660957f
C732 Vdd 17_8/a_26_538# 3.76551f
C733 GND 17_8/DATA 0.100362p
C734 17_23/a_252_786# 17_23/DATA 3.00456f
C735 GND 17_12/a_62_902# 2.79216f
C736 Vdd 17_17/DATA 0.111498p
C737 GND 17_15/OEN 4.46481f
C738 Vdd 17_15/DO 3.11769f
C739 GND 17_8/DI 4.11066f
C740 Vdd 17_12/DIB 6.39135f
C741 GND 17_12/a_58_538# 3.79746f
C742 Vdd 17_17/DI 3.31488f
C743 GND 17_17/a_62_82# 48.660957f
C744 GND 17_31/a_62_902# 2.79216f
C745 17_6/w_40_1480# p_c 66.6688f
C746 Vdd 17_31/DIB 6.39135f
C747 GND 17_31/a_58_538# 3.79746f
C748 Vdd 17_0/DO 3.11769f
C749 GND p_h 0.100362p
C750 Vdd 17_7/a_26_538# 3.79359f
C751 Vdd 17_27/DATA 0.111498p
C752 GND 17_25/OEN 4.46481f
C753 Vdd 17_25/DO 3.11769f
C754 GND 17_7/DI 4.11066f
C755 Vdd 17_27/DI 3.31488f
C756 GND 17_27/a_62_82# 48.660957f
C757 GND 17_35/OEN 4.46481f
C758 Vdd 17_35/DO 3.11769f
C759 17_6/a_420_786# p_c 2.95776f
C760 GND 17_20/a_62_902# 2.79216f
C761 17_9/a_62_902# 17_9/DATA 6.99264f
C762 Vdd 17_20/DIB 6.39135f
C763 GND 17_20/a_58_538# 3.79746f
C764 p_c 17_6/a_62_82# 8.056081f
C765 17_16/a_62_902# 17_16/DATA 6.99264f
C766 GND 17_1/OEN 4.46481f
C767 Vdd 17_1/DO 3.11769f
C768 17_11/a_62_902# 17_11/DATA 6.99264f
C769 Vdd 17_6/a_26_538# 3.76551f
C770 GND p_c 0.100362p
C771 17_13/a_252_786# 17_13/DATA 3.00456f
C772 Vdd 17_16/DATA 0.111498p
C773 GND 17_32/a_26_538# 3.75903f
C774 Vdd 17_16/DI 3.31488f
C775 GND 17_16/a_62_82# 48.660957f
C776 GND 17_34/OEN 4.46481f
C777 Vdd 17_34/DO 3.11769f
C778 GND 17_30/a_62_902# 2.79216f
C779 GND 17_32/m3_n72_n22# 32.52166f
C780 Vdd i 4.69701f
C781 17_5/w_40_1480# p_d 66.6688f
C782 Vdd 17_30/DIB 6.39135f
C783 GND 17_30/a_58_538# 3.79746f
C784 Vdd 17_5/a_26_538# 3.76551f
C785 GND p_d 0.100362p
C786 Vdd 17_26/DATA 0.111498p
C787 Vdd 18_0/w_40_1480# 66.6688f
C788 GND 17_21/a_26_538# 3.75903f
C789 17_35/m3_n72_n22# 0 5.6667f
C790 17_35/DI 0 28.906801f **FLOATING
C791 17_35/a_62_82# 0 49.1105f **FLOATING
C792 17_35/DIB 0 34.368f **FLOATING
C793 17_35/a_58_538# 0 8.3028f **FLOATING
C794 17_35/DO 0 15.5424f **FLOATING
C795 17_35/OEN 0 15.477599f **FLOATING
C796 17_35/a_26_538# 0 14.0407f **FLOATING
C797 17_35/DATA 0 0.227199p **FLOATING
C798 17_35/a_420_786# 0 5.0688f **FLOATING
C799 17_35/a_252_786# 0 5.148f **FLOATING
C800 17_35/a_62_902# 0 51.1622f **FLOATING
C801 17_35/w_40_1480# 0 0.237276p
C802 17_34/m3_n72_n22# 0 5.6667f
C803 17_34/DI 0 28.906801f **FLOATING
C804 17_34/a_62_82# 0 49.1105f **FLOATING
C805 17_34/DIB 0 34.368f **FLOATING
C806 17_34/a_58_538# 0 8.3028f **FLOATING
C807 17_34/DO 0 15.5424f **FLOATING
C808 17_34/OEN 0 15.477599f **FLOATING
C809 17_34/a_26_538# 0 14.0407f **FLOATING
C810 17_34/DATA 0 0.227199p **FLOATING
C811 17_34/a_420_786# 0 5.0688f **FLOATING
C812 17_34/a_252_786# 0 5.148f **FLOATING
C813 17_34/a_62_902# 0 51.1622f **FLOATING
C814 17_34/w_40_1480# 0 0.237276p
C815 17_24/m3_n72_n22# 0 5.6667f
C816 17_24/DI 0 28.906801f **FLOATING
C817 17_24/a_62_82# 0 49.1105f **FLOATING
C818 17_24/DIB 0 34.368f **FLOATING
C819 17_24/a_58_538# 0 8.3028f **FLOATING
C820 17_24/DO 0 15.5424f **FLOATING
C821 17_24/OEN 0 15.477599f **FLOATING
C822 17_24/a_26_538# 0 14.0407f **FLOATING
C823 17_24/DATA 0 0.227199p **FLOATING
C824 17_24/a_420_786# 0 5.0688f **FLOATING
C825 17_24/a_252_786# 0 5.148f **FLOATING
C826 17_24/a_62_902# 0 51.1622f **FLOATING
C827 17_24/w_40_1480# 0 0.237276p
C828 17_23/m3_n72_n22# 0 5.6667f
C829 17_23/DI 0 28.906801f **FLOATING
C830 17_23/a_62_82# 0 49.1105f **FLOATING
C831 17_23/DIB 0 34.368f **FLOATING
C832 17_23/a_58_538# 0 8.3028f **FLOATING
C833 17_23/DO 0 15.5424f **FLOATING
C834 17_23/OEN 0 15.477599f **FLOATING
C835 17_23/a_26_538# 0 14.0407f **FLOATING
C836 17_23/DATA 0 0.227199p **FLOATING
C837 17_23/a_420_786# 0 5.0688f **FLOATING
C838 17_23/a_252_786# 0 5.148f **FLOATING
C839 17_23/a_62_902# 0 51.1622f **FLOATING
C840 17_23/w_40_1480# 0 0.237276p
C841 17_13/m3_n72_n22# 0 5.6667f
C842 17_13/DI 0 28.906801f **FLOATING
C843 17_13/a_62_82# 0 49.1105f **FLOATING
C844 17_13/DIB 0 34.368f **FLOATING
C845 17_13/a_58_538# 0 8.3028f **FLOATING
C846 17_13/DO 0 15.5424f **FLOATING
C847 17_13/OEN 0 15.477599f **FLOATING
C848 17_13/a_26_538# 0 14.0407f **FLOATING
C849 17_13/DATA 0 0.227199p **FLOATING
C850 17_13/a_420_786# 0 5.0688f **FLOATING
C851 17_13/a_252_786# 0 5.148f **FLOATING
C852 17_13/a_62_902# 0 51.1622f **FLOATING
C853 17_13/w_40_1480# 0 0.237276p
C854 17_12/m3_n72_n22# 0 5.6667f
C855 17_12/DI 0 28.906801f **FLOATING
C856 17_12/a_62_82# 0 49.1105f **FLOATING
C857 17_12/DIB 0 34.368f **FLOATING
C858 17_12/a_58_538# 0 8.3028f **FLOATING
C859 17_12/DO 0 15.5424f **FLOATING
C860 17_12/OEN 0 15.477599f **FLOATING
C861 17_12/a_26_538# 0 14.0407f **FLOATING
C862 17_12/DATA 0 0.227199p **FLOATING
C863 17_12/a_420_786# 0 5.0688f **FLOATING
C864 17_12/a_252_786# 0 5.148f **FLOATING
C865 17_12/a_62_902# 0 51.1622f **FLOATING
C866 17_12/w_40_1480# 0 0.237276p
C867 17_33/m3_n72_n22# 0 5.6667f
C868 17_33/DI 0 28.906801f **FLOATING
C869 17_33/a_62_82# 0 49.1105f **FLOATING
C870 17_33/DIB 0 34.368f **FLOATING
C871 17_33/a_58_538# 0 8.3028f **FLOATING
C872 17_33/DO 0 15.5424f **FLOATING
C873 17_33/OEN 0 15.477599f **FLOATING
C874 17_33/a_26_538# 0 14.0407f **FLOATING
C875 17_33/DATA 0 0.227199p **FLOATING
C876 17_33/a_420_786# 0 5.0688f **FLOATING
C877 17_33/a_252_786# 0 5.148f **FLOATING
C878 17_33/a_62_902# 0 51.1622f **FLOATING
C879 17_33/w_40_1480# 0 0.237276p
C880 17_22/m3_n72_n22# 0 5.6667f
C881 17_22/DI 0 28.906801f **FLOATING
C882 17_22/a_62_82# 0 49.1105f **FLOATING
C883 17_22/DIB 0 34.368f **FLOATING
C884 17_22/a_58_538# 0 8.3028f **FLOATING
C885 17_22/DO 0 15.5424f **FLOATING
C886 17_22/OEN 0 15.477599f **FLOATING
C887 17_22/a_26_538# 0 14.0407f **FLOATING
C888 17_22/DATA 0 0.227199p **FLOATING
C889 17_22/a_420_786# 0 5.0688f **FLOATING
C890 17_22/a_252_786# 0 5.148f **FLOATING
C891 17_22/a_62_902# 0 51.1622f **FLOATING
C892 17_22/w_40_1480# 0 0.237276p
C893 17_11/m3_n72_n22# 0 5.6667f
C894 17_11/DI 0 28.906801f **FLOATING
C895 17_11/a_62_82# 0 49.1105f **FLOATING
C896 17_11/DIB 0 34.368f **FLOATING
C897 17_11/a_58_538# 0 8.3028f **FLOATING
C898 17_11/DO 0 15.5424f **FLOATING
C899 17_11/OEN 0 15.477599f **FLOATING
C900 17_11/a_26_538# 0 14.0407f **FLOATING
C901 17_11/DATA 0 0.227199p **FLOATING
C902 17_11/a_420_786# 0 5.0688f **FLOATING
C903 17_11/a_252_786# 0 5.148f **FLOATING
C904 17_11/a_62_902# 0 51.1622f **FLOATING
C905 17_11/w_40_1480# 0 0.237276p
C906 17_32/m3_n72_n22# 0 5.6667f
C907 17_32/DI 0 28.906801f **FLOATING
C908 17_32/a_62_82# 0 49.1105f **FLOATING
C909 17_32/DIB 0 34.368f **FLOATING
C910 17_32/a_58_538# 0 8.3028f **FLOATING
C911 17_32/DO 0 15.5424f **FLOATING
C912 17_32/OEN 0 15.477599f **FLOATING
C913 17_32/a_26_538# 0 14.0407f **FLOATING
C914 17_32/DATA 0 0.227199p **FLOATING
C915 17_32/a_420_786# 0 5.0688f **FLOATING
C916 17_32/a_252_786# 0 5.148f **FLOATING
C917 17_32/a_62_902# 0 51.1622f **FLOATING
C918 17_32/w_40_1480# 0 0.237276p
C919 17_21/m3_n72_n22# 0 5.6667f
C920 17_21/DI 0 28.906801f **FLOATING
C921 17_21/a_62_82# 0 49.1105f **FLOATING
C922 17_21/DIB 0 34.368f **FLOATING
C923 17_21/a_58_538# 0 8.3028f **FLOATING
C924 17_21/DO 0 15.5424f **FLOATING
C925 17_21/OEN 0 15.477599f **FLOATING
C926 17_21/a_26_538# 0 14.0407f **FLOATING
C927 17_21/DATA 0 0.227199p **FLOATING
C928 17_21/a_420_786# 0 5.0688f **FLOATING
C929 17_21/a_252_786# 0 5.148f **FLOATING
C930 17_21/a_62_902# 0 51.1622f **FLOATING
C931 17_21/w_40_1480# 0 0.237276p
C932 17_10/m3_n72_n22# 0 5.6667f
C933 17_10/DI 0 28.906801f **FLOATING
C934 17_10/a_62_82# 0 49.1105f **FLOATING
C935 17_10/DIB 0 34.368f **FLOATING
C936 17_10/a_58_538# 0 8.3028f **FLOATING
C937 17_10/DO 0 15.5424f **FLOATING
C938 17_10/OEN 0 15.477599f **FLOATING
C939 17_10/a_26_538# 0 14.0407f **FLOATING
C940 17_10/DATA 0 0.227199p **FLOATING
C941 17_10/a_420_786# 0 5.0688f **FLOATING
C942 17_10/a_252_786# 0 5.148f **FLOATING
C943 17_10/a_62_902# 0 51.1622f **FLOATING
C944 17_10/w_40_1480# 0 0.237276p
C945 18_1/w_40_1480# 0 0.237276p
C946 17_31/m3_n72_n22# 0 5.6667f
C947 17_31/DI 0 28.906801f **FLOATING
C948 17_31/a_62_82# 0 49.1105f **FLOATING
C949 17_31/DIB 0 34.368f **FLOATING
C950 17_31/a_58_538# 0 8.3028f **FLOATING
C951 17_31/DO 0 15.5424f **FLOATING
C952 17_31/OEN 0 15.477599f **FLOATING
C953 17_31/a_26_538# 0 14.0407f **FLOATING
C954 17_31/DATA 0 0.227199p **FLOATING
C955 17_31/a_420_786# 0 5.0688f **FLOATING
C956 17_31/a_252_786# 0 5.148f **FLOATING
C957 17_31/a_62_902# 0 51.1622f **FLOATING
C958 17_31/w_40_1480# 0 0.237276p
C959 17_20/m3_n72_n22# 0 5.6667f
C960 17_20/DI 0 28.906801f **FLOATING
C961 17_20/a_62_82# 0 49.1105f **FLOATING
C962 17_20/DIB 0 34.368f **FLOATING
C963 17_20/a_58_538# 0 8.3028f **FLOATING
C964 17_20/DO 0 15.5424f **FLOATING
C965 17_20/OEN 0 15.477599f **FLOATING
C966 17_20/a_26_538# 0 14.0407f **FLOATING
C967 17_20/DATA 0 0.227199p **FLOATING
C968 17_20/a_420_786# 0 5.0688f **FLOATING
C969 17_20/a_252_786# 0 5.148f **FLOATING
C970 17_20/a_62_902# 0 51.1622f **FLOATING
C971 17_20/w_40_1480# 0 0.237276p
C972 17_30/m3_n72_n22# 0 5.6667f
C973 17_30/DI 0 28.906801f **FLOATING
C974 17_30/a_62_82# 0 49.1105f **FLOATING
C975 17_30/DIB 0 34.368f **FLOATING
C976 17_30/a_58_538# 0 8.3028f **FLOATING
C977 17_30/DO 0 15.5424f **FLOATING
C978 17_30/OEN 0 15.477599f **FLOATING
C979 17_30/a_26_538# 0 14.0407f **FLOATING
C980 17_30/DATA 0 0.227199p **FLOATING
C981 17_30/a_420_786# 0 5.0688f **FLOATING
C982 17_30/a_252_786# 0 5.148f **FLOATING
C983 17_30/a_62_902# 0 51.1622f **FLOATING
C984 17_30/w_40_1480# 0 0.237276p
C985 18_0/w_40_1480# 0 0.237276p
C986 17_9/m3_n72_n22# 0 5.6667f
C987 17_9/DI 0 28.906801f **FLOATING
C988 17_9/a_62_82# 0 49.1105f **FLOATING
C989 17_9/DIB 0 34.368f **FLOATING
C990 17_9/a_58_538# 0 8.3028f **FLOATING
C991 17_9/DO 0 15.5424f **FLOATING
C992 17_9/OEN 0 15.477599f **FLOATING
C993 17_9/a_26_538# 0 14.0407f **FLOATING
C994 17_9/DATA 0 0.227199p **FLOATING
C995 17_9/a_420_786# 0 5.0688f **FLOATING
C996 17_9/a_252_786# 0 5.148f **FLOATING
C997 17_9/a_62_902# 0 51.1622f **FLOATING
C998 17_9/w_40_1480# 0 0.237276p
C999 17_8/m3_n72_n22# 0 5.6667f
C1000 17_8/DI 0 28.906801f **FLOATING
C1001 17_8/a_62_82# 0 49.1105f **FLOATING
C1002 17_8/DIB 0 34.368f **FLOATING
C1003 17_8/a_58_538# 0 8.3028f **FLOATING
C1004 17_8/DO 0 15.5424f **FLOATING
C1005 17_8/OEN 0 15.477599f **FLOATING
C1006 17_8/a_26_538# 0 14.0407f **FLOATING
C1007 17_8/DATA 0 0.227199p **FLOATING
C1008 17_8/a_420_786# 0 5.0688f **FLOATING
C1009 17_8/a_252_786# 0 5.148f **FLOATING
C1010 17_8/a_62_902# 0 51.1622f **FLOATING
C1011 17_8/w_40_1480# 0 0.237276p
C1012 17_7/m3_n72_n22# 0 5.6667f
C1013 17_7/DI 0 28.906801f **FLOATING
C1014 17_7/a_62_82# 0 49.1105f **FLOATING
C1015 17_7/DIB 0 34.368f **FLOATING
C1016 17_7/a_58_538# 0 8.3028f **FLOATING
C1017 17_7/a_26_538# 0 14.0407f **FLOATING
C1018 p_h 0 0.222516p **FLOATING
C1019 17_7/a_420_786# 0 5.0688f **FLOATING
C1020 17_7/a_252_786# 0 5.148f **FLOATING
C1021 17_7/a_62_902# 0 51.1622f **FLOATING
C1022 17_7/w_40_1480# 0 0.237276p
C1023 17_6/m3_n72_n22# 0 5.6667f
C1024 17_6/a_62_82# 0 49.1105f **FLOATING
C1025 17_6/DIB 0 34.368f **FLOATING
C1026 17_6/a_58_538# 0 8.3028f **FLOATING
C1027 17_6/DO 0 15.5424f **FLOATING
C1028 17_6/a_26_538# 0 14.0407f **FLOATING
C1029 p_c 0 0.2228p **FLOATING
C1030 17_6/a_420_786# 0 5.0688f **FLOATING
C1031 17_6/a_252_786# 0 5.148f **FLOATING
C1032 17_6/a_62_902# 0 51.1622f **FLOATING
C1033 17_6/w_40_1480# 0 0.237276p
C1034 17_5/m3_n72_n22# 0 5.6667f
C1035 17_5/a_62_82# 0 49.1105f **FLOATING
C1036 17_5/DIB 0 34.368f **FLOATING
C1037 17_5/a_58_538# 0 8.3028f **FLOATING
C1038 17_5/DO 0 15.5424f **FLOATING
C1039 17_5/a_26_538# 0 14.0407f **FLOATING
C1040 p_d 0 0.221663p **FLOATING
C1041 17_5/a_420_786# 0 5.0688f **FLOATING
C1042 17_5/a_252_786# 0 5.148f **FLOATING
C1043 17_5/a_62_902# 0 51.1622f **FLOATING
C1044 17_5/w_40_1480# 0 0.237276p
C1045 17_4/m3_n72_n22# 0 5.6667f
C1046 17_4/a_62_82# 0 49.1105f **FLOATING
C1047 17_4/DIB 0 34.368f **FLOATING
C1048 17_4/a_58_538# 0 8.3028f **FLOATING
C1049 17_4/DO 0 15.5424f **FLOATING
C1050 17_4/a_26_538# 0 14.0407f **FLOATING
C1051 p_b 0 0.223673p **FLOATING
C1052 17_4/a_420_786# 0 5.0688f **FLOATING
C1053 17_4/a_252_786# 0 5.148f **FLOATING
C1054 17_4/a_62_902# 0 51.1622f **FLOATING
C1055 17_4/w_40_1480# 0 0.237276p
C1056 17_3/m3_n72_n22# 0 5.6667f
C1057 17_3/DI 0 28.906801f **FLOATING
C1058 17_3/a_62_82# 0 49.1105f **FLOATING
C1059 17_3/DIB 0 34.368f **FLOATING
C1060 17_3/a_58_538# 0 8.3028f **FLOATING
C1061 17_3/a_26_538# 0 14.0407f **FLOATING
C1062 p_i 0 0.227199p **FLOATING
C1063 17_3/a_420_786# 0 5.0688f **FLOATING
C1064 17_3/a_252_786# 0 5.148f **FLOATING
C1065 17_3/a_62_902# 0 51.1622f **FLOATING
C1066 17_3/w_40_1480# 0 0.237276p
C1067 17_2/m3_n72_n22# 0 5.6667f
C1068 17_2/a_62_82# 0 49.1105f **FLOATING
C1069 17_2/DIB 0 34.368f **FLOATING
C1070 17_2/a_58_538# 0 8.3028f **FLOATING
C1071 17_2/DO 0 15.5424f **FLOATING
C1072 17_2/a_26_538# 0 14.0407f **FLOATING
C1073 p_a 0 0.220953p **FLOATING
C1074 17_2/a_420_786# 0 5.0688f **FLOATING
C1075 17_2/a_252_786# 0 5.148f **FLOATING
C1076 17_2/a_62_902# 0 51.1622f **FLOATING
C1077 17_2/w_40_1480# 0 0.237276p
C1078 17_0/m3_n72_n22# 0 5.6667f
C1079 17_0/DI 0 28.906801f **FLOATING
C1080 17_0/a_62_82# 0 49.1105f **FLOATING
C1081 17_0/DIB 0 34.368f **FLOATING
C1082 17_0/a_58_538# 0 8.3028f **FLOATING
C1083 17_0/DO 0 15.5424f **FLOATING
C1084 17_0/a_26_538# 0 14.0407f **FLOATING
C1085 17_0/DATA 0 0.227199p **FLOATING
C1086 17_0/a_420_786# 0 5.0688f **FLOATING
C1087 17_0/a_252_786# 0 5.148f **FLOATING
C1088 17_0/a_62_902# 0 51.1622f **FLOATING
C1089 17_0/w_40_1480# 0 0.237276p
C1090 17_1/m3_n72_n22# 0 5.6667f
C1091 17_1/DI 0 28.906801f **FLOATING
C1092 17_1/a_62_82# 0 49.1105f **FLOATING
C1093 17_1/DIB 0 34.368f **FLOATING
C1094 17_1/a_58_538# 0 8.3028f **FLOATING
C1095 17_1/DO 0 15.5424f **FLOATING
C1096 17_1/OEN 0 15.477599f **FLOATING
C1097 17_1/a_26_538# 0 14.0407f **FLOATING
C1098 17_1/DATA 0 0.227199p **FLOATING
C1099 17_1/a_420_786# 0 5.0688f **FLOATING
C1100 17_1/a_252_786# 0 5.148f **FLOATING
C1101 17_1/a_62_902# 0 51.1622f **FLOATING
C1102 17_1/w_40_1480# 0 0.237276p
C1103 19_1/w_40_1480# 0 0.237276p
C1104 19_0/w_40_1480# 0 0.237276p
C1105 17_19/m3_n72_n22# 0 5.6667f
C1106 17_19/DI 0 28.906801f **FLOATING
C1107 17_19/a_62_82# 0 49.1105f **FLOATING
C1108 17_19/DIB 0 34.368f **FLOATING
C1109 17_19/a_58_538# 0 8.3028f **FLOATING
C1110 17_19/DO 0 15.5424f **FLOATING
C1111 17_19/OEN 0 15.477599f **FLOATING
C1112 17_19/a_26_538# 0 14.0407f **FLOATING
C1113 17_19/DATA 0 0.227199p **FLOATING
C1114 17_19/a_420_786# 0 5.0688f **FLOATING
C1115 17_19/a_252_786# 0 5.148f **FLOATING
C1116 17_19/a_62_902# 0 51.1622f **FLOATING
C1117 17_19/w_40_1480# 0 0.237276p
C1118 17_29/m3_n72_n22# 0 5.6667f
C1119 17_29/DI 0 28.906801f **FLOATING
C1120 17_29/a_62_82# 0 49.1105f **FLOATING
C1121 17_29/DIB 0 34.368f **FLOATING
C1122 17_29/a_58_538# 0 8.3028f **FLOATING
C1123 17_29/DO 0 15.5424f **FLOATING
C1124 17_29/OEN 0 15.477599f **FLOATING
C1125 17_29/a_26_538# 0 14.0407f **FLOATING
C1126 17_29/DATA 0 0.227199p **FLOATING
C1127 17_29/a_420_786# 0 5.0688f **FLOATING
C1128 17_29/a_252_786# 0 5.148f **FLOATING
C1129 17_29/a_62_902# 0 51.1622f **FLOATING
C1130 17_29/w_40_1480# 0 0.237276p
C1131 h 0 0.309389p **FLOATING
C1132 hwtest_0/AND2X2_0/a_4_12# 0 6.03567f **FLOATING
C1133 c 0 0.166913p **FLOATING
C1134 hwtest_0/NOR2X1_1/Y 0 6.23106f **FLOATING
C1135 d 0 0.136841p **FLOATING
C1136 i 0 0.316458p **FLOATING
C1137 a 0 0.25947p **FLOATING
C1138 b 0 0.211135p **FLOATING
C1139 17_18/m3_n72_n22# 0 5.6667f
C1140 17_18/DI 0 28.906801f **FLOATING
C1141 17_18/a_62_82# 0 49.1105f **FLOATING
C1142 17_18/DIB 0 34.368f **FLOATING
C1143 17_18/a_58_538# 0 8.3028f **FLOATING
C1144 17_18/DO 0 15.5424f **FLOATING
C1145 17_18/OEN 0 15.477599f **FLOATING
C1146 17_18/a_26_538# 0 14.0407f **FLOATING
C1147 17_18/DATA 0 0.227199p **FLOATING
C1148 17_18/a_420_786# 0 5.0688f **FLOATING
C1149 17_18/a_252_786# 0 5.148f **FLOATING
C1150 17_18/a_62_902# 0 51.1622f **FLOATING
C1151 17_18/w_40_1480# 0 0.237276p
C1152 17_28/m3_n72_n22# 0 5.6667f
C1153 17_28/DI 0 28.906801f **FLOATING
C1154 17_28/a_62_82# 0 49.1105f **FLOATING
C1155 17_28/DIB 0 34.368f **FLOATING
C1156 17_28/a_58_538# 0 8.3028f **FLOATING
C1157 17_28/DO 0 15.5424f **FLOATING
C1158 17_28/OEN 0 15.477599f **FLOATING
C1159 17_28/a_26_538# 0 14.0407f **FLOATING
C1160 17_28/DATA 0 0.227199p **FLOATING
C1161 17_28/a_420_786# 0 5.0688f **FLOATING
C1162 17_28/a_252_786# 0 5.148f **FLOATING
C1163 17_28/a_62_902# 0 51.1622f **FLOATING
C1164 17_28/w_40_1480# 0 0.237276p
C1165 17_17/m3_n72_n22# 0 5.6667f
C1166 17_17/DI 0 28.906801f **FLOATING
C1167 17_17/a_62_82# 0 49.1105f **FLOATING
C1168 17_17/DIB 0 34.368f **FLOATING
C1169 17_17/a_58_538# 0 8.3028f **FLOATING
C1170 17_17/DO 0 15.5424f **FLOATING
C1171 17_17/OEN 0 15.477599f **FLOATING
C1172 17_17/a_26_538# 0 14.0407f **FLOATING
C1173 17_17/DATA 0 0.227199p **FLOATING
C1174 17_17/a_420_786# 0 5.0688f **FLOATING
C1175 17_17/a_252_786# 0 5.148f **FLOATING
C1176 17_17/a_62_902# 0 51.1622f **FLOATING
C1177 17_17/w_40_1480# 0 0.237276p
C1178 17_27/m3_n72_n22# 0 5.6667f
C1179 17_27/DI 0 28.906801f **FLOATING
C1180 17_27/a_62_82# 0 49.1105f **FLOATING
C1181 17_27/DIB 0 34.368f **FLOATING
C1182 17_27/a_58_538# 0 8.3028f **FLOATING
C1183 17_27/DO 0 15.5424f **FLOATING
C1184 17_27/OEN 0 15.477599f **FLOATING
C1185 17_27/a_26_538# 0 14.0407f **FLOATING
C1186 17_27/DATA 0 0.227199p **FLOATING
C1187 17_27/a_420_786# 0 5.0688f **FLOATING
C1188 17_27/a_252_786# 0 5.148f **FLOATING
C1189 17_27/a_62_902# 0 51.1622f **FLOATING
C1190 17_27/w_40_1480# 0 0.237276p
C1191 17_16/m3_n72_n22# 0 5.6667f
C1192 17_16/DI 0 28.906801f **FLOATING
C1193 17_16/a_62_82# 0 49.1105f **FLOATING
C1194 17_16/DIB 0 34.368f **FLOATING
C1195 17_16/a_58_538# 0 8.3028f **FLOATING
C1196 17_16/DO 0 15.5424f **FLOATING
C1197 17_16/OEN 0 15.477599f **FLOATING
C1198 17_16/a_26_538# 0 14.0407f **FLOATING
C1199 17_16/DATA 0 0.227199p **FLOATING
C1200 17_16/a_420_786# 0 5.0688f **FLOATING
C1201 17_16/a_252_786# 0 5.148f **FLOATING
C1202 17_16/a_62_902# 0 51.1622f **FLOATING
C1203 17_16/w_40_1480# 0 0.237276p
C1204 17_26/DI 0 28.906801f **FLOATING
C1205 17_26/a_62_82# 0 49.1105f **FLOATING
C1206 17_26/DIB 0 34.368f **FLOATING
C1207 17_26/a_58_538# 0 8.3028f **FLOATING
C1208 17_26/DO 0 15.5424f **FLOATING
C1209 17_26/OEN 0 15.477599f **FLOATING
C1210 17_26/a_26_538# 0 14.0407f **FLOATING
C1211 17_26/DATA 0 0.227199p **FLOATING
C1212 17_26/a_420_786# 0 5.0688f **FLOATING
C1213 17_26/a_252_786# 0 5.148f **FLOATING
C1214 17_26/a_62_902# 0 51.1622f **FLOATING
C1215 17_26/w_40_1480# 0 0.237276p
C1216 17_15/m3_n72_n22# 0 5.6667f
C1217 17_15/DI 0 28.906801f **FLOATING
C1218 17_15/a_62_82# 0 49.1105f **FLOATING
C1219 17_15/DIB 0 34.368f **FLOATING
C1220 17_15/a_58_538# 0 8.3028f **FLOATING
C1221 17_15/DO 0 15.5424f **FLOATING
C1222 17_15/OEN 0 15.477599f **FLOATING
C1223 17_15/a_26_538# 0 14.0407f **FLOATING
C1224 17_15/DATA 0 0.227199p **FLOATING
C1225 17_15/a_420_786# 0 5.0688f **FLOATING
C1226 17_15/a_252_786# 0 5.148f **FLOATING
C1227 17_15/a_62_902# 0 51.1622f **FLOATING
C1228 17_15/w_40_1480# 0 0.237276p
C1229 17_26/m3_n72_n22# 0 9.5652f
C1230 17_25/DI 0 28.906801f **FLOATING
C1231 17_25/a_62_82# 0 49.1105f **FLOATING
C1232 17_25/DIB 0 34.368f **FLOATING
C1233 17_25/a_58_538# 0 8.3028f **FLOATING
C1234 17_25/DO 0 15.5424f **FLOATING
C1235 17_25/OEN 0 15.477599f **FLOATING
C1236 17_25/a_26_538# 0 14.0407f **FLOATING
C1237 17_25/DATA 0 0.227199p **FLOATING
C1238 17_25/a_420_786# 0 5.0688f **FLOATING
C1239 17_25/a_252_786# 0 5.148f **FLOATING
C1240 17_25/a_62_902# 0 51.1622f **FLOATING
C1241 17_25/w_40_1480# 0 0.237276p
C1242 Vdd 0 20.958416p **FLOATING
C1243 17_14/m3_n72_n22# 0 5.6667f
C1244 17_14/DI 0 28.906801f **FLOATING
C1245 17_14/a_62_82# 0 49.1105f **FLOATING
C1246 17_14/DIB 0 34.368f **FLOATING
C1247 17_14/a_58_538# 0 8.3028f **FLOATING
C1248 17_14/DO 0 15.5424f **FLOATING
C1249 17_14/OEN 0 15.477599f **FLOATING
C1250 17_14/a_26_538# 0 14.0407f **FLOATING
C1251 17_14/DATA 0 0.227199p **FLOATING
C1252 17_14/a_420_786# 0 5.0688f **FLOATING
C1253 17_14/a_252_786# 0 5.148f **FLOATING
C1254 17_14/a_62_902# 0 51.1622f **FLOATING
C1255 17_14/w_40_1480# 0 0.237276p
