magic
tech scmos
timestamp 1712112060
<< end >>
