magic
tech scmos
timestamp 1714524305
<< m2contact >>
rect -2 -2 2 2
<< end >>
