magic
tech scmos
timestamp 1712111715
<< end >>
