magic
tech scmos
timestamp 1714528750
<< nwell >>
rect -1158 1473 -1141 1485
rect -858 1470 -837 1486
rect -560 1468 -545 1484
rect -1090 1449 -1077 1465
rect -792 1447 -777 1462
rect -491 1450 -477 1464
rect 1478 1457 1490 1470
rect -1446 1218 -1433 1230
rect 1466 1157 1478 1170
rect -406 1048 -391 1077
rect -327 1058 -282 1094
rect -232 1069 -187 1105
rect -1331 945 -1316 957
rect -1454 921 -1441 933
rect 1365 856 1391 883
rect 1408 549 1430 565
rect -1285 531 -1270 543
rect -1403 427 -1382 440
rect -1318 363 -1282 384
rect 1455 248 1471 266
rect -1224 -245 -1197 -227
rect -1426 -343 -1411 -329
rect -1182 -340 -1155 -322
rect 1361 -344 1388 -328
rect 321 -1436 333 -1422
rect 394 -1435 406 -1421
<< metal1 >>
rect -1156 1485 -1147 1489
rect -1155 1418 -1147 1473
rect -1090 1465 -1085 1490
rect -864 1486 -846 1487
rect -864 1470 -858 1486
rect -1490 1311 -1409 1317
rect -1444 1289 -1434 1311
rect -1446 1230 -1434 1289
rect -1310 1244 -1285 1252
rect -1161 1071 -1140 1418
rect -864 1404 -846 1470
rect -792 1462 -777 1495
rect -559 1484 -544 1489
rect -545 1468 -544 1484
rect -493 1485 -480 1491
rect -493 1474 -478 1485
rect -867 1153 -846 1404
rect -559 1340 -544 1468
rect -491 1464 -478 1474
rect 1452 1457 1478 1466
rect 1253 1416 1336 1422
rect 1452 1416 1463 1457
rect 1253 1386 1463 1416
rect -568 1220 -536 1340
rect 1253 1248 1336 1386
rect 1229 1239 1336 1248
rect -222 1220 -194 1225
rect -568 1196 -182 1220
rect -867 1115 -296 1153
rect -866 1112 -296 1115
rect -325 1094 -298 1112
rect -222 1105 -194 1196
rect -1161 1048 -406 1071
rect -1161 1042 -391 1048
rect -1161 1039 -1140 1042
rect -1491 1011 -1430 1017
rect -1452 992 -1440 1011
rect -1454 983 -1440 992
rect -1454 933 -1441 983
rect -1332 957 -1314 1006
rect 1155 992 1197 997
rect 1229 992 1276 1239
rect -1332 945 -1331 957
rect -1316 945 -1314 957
rect 1154 959 1276 992
rect 1305 1167 1347 1175
rect 1305 1157 1466 1167
rect 1478 1166 1479 1167
rect 1478 1157 1487 1166
rect 1305 1154 1462 1157
rect 1154 955 1266 959
rect -1332 790 -1314 945
rect -1333 780 -1314 790
rect -1333 578 -1315 780
rect 1155 614 1197 955
rect 1305 618 1347 1154
rect 1362 856 1365 864
rect 973 579 1255 614
rect 1155 578 1197 579
rect -1333 564 -1231 578
rect 1305 531 1345 618
rect 1078 482 1345 531
rect 1362 466 1390 856
rect 1404 565 1437 566
rect 1404 549 1408 565
rect 1430 549 1437 565
rect 1027 438 1392 466
rect -1382 427 -1290 437
rect 1362 436 1390 438
rect 1404 275 1437 549
rect -1426 245 -1305 256
rect 1132 245 1437 275
rect 1454 266 1470 267
rect 1454 258 1455 266
rect 1454 248 1455 254
rect -1425 60 -1411 245
rect 1132 243 1413 245
rect 1332 232 1433 233
rect 1454 232 1470 248
rect 1332 219 1474 232
rect 1332 67 1433 219
rect -1426 -329 -1411 60
rect 1360 -328 1386 46
rect 1360 -344 1361 -328
rect 1360 -357 1386 -344
rect -1405 -643 -1382 -620
rect -1343 -944 -1315 -930
rect -858 -1012 -792 -1007
rect -858 -1070 -855 -1012
rect -1297 -1255 -1252 -1217
rect -858 -1444 -792 -1070
rect 333 -1435 394 -1423
rect 333 -1436 402 -1435
rect -856 -1480 -841 -1444
rect -846 -1486 -841 -1480
rect -789 -1489 -784 -1470
<< m2contact >>
rect -1158 1473 -1141 1485
rect -858 1470 -837 1486
rect -1090 1449 -1077 1465
rect -1446 1218 -1433 1230
rect -560 1468 -545 1484
rect -792 1447 -777 1462
rect -491 1450 -477 1464
rect 1478 1457 1490 1470
rect -406 1048 -391 1077
rect -327 1058 -282 1094
rect -232 1069 -187 1105
rect -1454 921 -1441 933
rect -1331 945 -1316 957
rect 1466 1157 1478 1170
rect 1365 856 1391 883
rect -1285 531 -1270 543
rect 1408 549 1430 565
rect -1403 427 -1382 440
rect -1318 363 -1282 384
rect 1455 248 1471 266
rect -1224 -245 -1197 -227
rect -1426 -343 -1411 -329
rect -1182 -340 -1155 -322
rect 1361 -344 1388 -328
rect -855 -1070 -790 -1012
rect 340 -1340 376 -1301
rect 321 -1436 333 -1422
rect 394 -1435 406 -1421
rect -795 -1470 -784 -1462
rect -856 -1486 -846 -1480
<< metal2 >>
rect -1477 1476 -1471 1486
rect -1406 1476 -1400 1490
rect -1477 1470 -1400 1476
rect -1243 1412 -1234 1485
rect -1179 1463 -1170 1483
rect -1179 1462 -1106 1463
rect -1179 1450 -1090 1462
rect -1106 1449 -1090 1450
rect -878 1461 -869 1491
rect -878 1448 -792 1461
rect -878 1446 -869 1448
rect -862 1446 -818 1448
rect -777 1448 -772 1461
rect -578 1457 -570 1486
rect -506 1457 -491 1458
rect -578 1450 -491 1457
rect -277 1462 -272 1492
rect -206 1462 -201 1492
rect -477 1450 -471 1458
rect -578 1449 -502 1450
rect -578 1448 -570 1449
rect -277 1448 -197 1462
rect -42 1452 -35 1486
rect 21 1461 30 1486
rect 92 1461 99 1492
rect -276 1447 -197 1448
rect -1243 1407 -1233 1412
rect -1242 1353 -1233 1407
rect -1485 1244 -1283 1253
rect -1484 1230 -1429 1232
rect -1484 1222 -1446 1230
rect -1433 1222 -1429 1230
rect -1248 993 -1231 1353
rect -65 1106 -34 1452
rect 21 1451 100 1461
rect 257 1355 270 1486
rect 623 1447 629 1485
rect 692 1447 698 1495
rect 623 1437 702 1447
rect 692 1436 698 1437
rect 246 1347 303 1355
rect 70 1342 303 1347
rect 65 1312 303 1342
rect 65 1106 105 1312
rect 246 1311 303 1312
rect 257 1309 270 1311
rect 858 1273 876 1486
rect 922 1441 928 1483
rect 993 1441 998 1493
rect 922 1424 1011 1441
rect 993 1423 998 1424
rect 278 1270 880 1273
rect 273 1223 880 1270
rect 273 1114 293 1223
rect 1160 1207 1180 1487
rect 1224 1463 1229 1483
rect 1294 1463 1300 1489
rect 1223 1454 1307 1463
rect 1294 1453 1300 1454
rect 1458 1294 1495 1299
rect 1458 1230 1466 1294
rect 1458 1223 1487 1230
rect 1027 1121 1192 1207
rect 1462 1166 1466 1167
rect 1461 1157 1466 1166
rect 1478 1166 1479 1167
rect 1478 1157 1487 1166
rect 450 1071 1192 1121
rect 1027 1061 1192 1071
rect -1243 975 -1231 993
rect 1462 995 1492 999
rect -1248 969 -776 975
rect -1248 967 -737 969
rect -1484 945 -1331 953
rect -1316 945 -1315 953
rect -1243 951 -737 967
rect -1484 944 -1315 945
rect -1485 922 -1454 930
rect -1441 922 -1436 930
rect 1462 929 1474 995
rect 1462 922 1486 929
rect -1358 865 -1352 867
rect -1485 856 -1352 865
rect -1490 695 -1438 698
rect -1444 630 -1438 695
rect -1483 622 -1435 630
rect -1488 567 -1383 569
rect -1488 556 -1382 567
rect -1403 440 -1382 556
rect -1358 542 -1352 856
rect 1363 856 1365 867
rect 1391 858 1488 867
rect 1391 856 1474 858
rect 1363 855 1474 856
rect 1457 699 1471 701
rect 1457 694 1496 699
rect 1457 630 1471 694
rect 1457 624 1487 630
rect 1457 623 1471 624
rect 1404 565 1486 566
rect 1404 556 1408 565
rect 1430 556 1486 565
rect -1358 532 -1285 542
rect -1270 532 -1248 542
rect 1462 401 1474 402
rect -1492 395 -1462 400
rect -1471 329 -1462 395
rect 1462 394 1496 401
rect -1332 363 -1318 383
rect -1485 324 -1457 329
rect -1453 319 -1442 337
rect -1332 334 -1283 363
rect -1393 319 -1283 334
rect 1462 330 1474 394
rect 1462 323 1492 330
rect -1453 301 -1283 319
rect -1453 296 -1337 301
rect -1484 -29 -1465 -23
rect -1476 -93 -1466 -29
rect -1493 -100 -1466 -93
rect -1476 -101 -1466 -100
rect -1453 -257 -1442 296
rect 1471 258 1486 266
rect 1486 243 1491 254
rect 1466 99 1494 100
rect 1465 95 1494 99
rect 1465 29 1474 95
rect 1465 21 1483 29
rect -1225 -245 -1224 -227
rect -1485 -266 -1412 -257
rect -1487 -343 -1426 -329
rect -1411 -343 -1410 -329
rect -1489 -505 -1451 -501
rect -1464 -570 -1452 -505
rect -1486 -577 -1452 -570
rect -1405 -632 -1382 -620
rect -1487 -643 -1382 -632
rect -1459 -800 -1453 -799
rect -1491 -805 -1453 -800
rect -1459 -870 -1453 -805
rect -1485 -875 -1448 -870
rect -1459 -877 -1453 -875
rect -1343 -934 -1315 -930
rect -1485 -944 -1315 -934
rect -1488 -1105 -1432 -1098
rect -1443 -1173 -1434 -1105
rect -1486 -1180 -1430 -1173
rect -1225 -1206 -1199 -245
rect -1297 -1230 -1252 -1217
rect -1486 -1244 -1252 -1230
rect -1297 -1255 -1252 -1244
rect -1236 -1223 -1199 -1206
rect -1184 -322 -1158 -308
rect -1184 -340 -1182 -322
rect -1470 -1400 -1456 -1394
rect -1236 -1399 -1209 -1223
rect -1184 -1277 -1158 -340
rect 1388 -344 1491 -334
rect 1465 -501 1495 -500
rect 1464 -506 1495 -501
rect 1464 -570 1474 -506
rect 1464 -577 1488 -570
rect -1184 -1299 -924 -1277
rect -1184 -1304 -1158 -1299
rect -1492 -1404 -1456 -1400
rect -1470 -1466 -1456 -1404
rect -1243 -1406 -1209 -1399
rect -1476 -1469 -1390 -1466
rect -1484 -1476 -1390 -1469
rect -1476 -1486 -1463 -1476
rect -1405 -1491 -1398 -1476
rect -1243 -1486 -1225 -1406
rect -1177 -1474 -1097 -1469
rect -1177 -1485 -1169 -1474
rect -1105 -1489 -1099 -1474
rect -942 -1485 -929 -1299
rect -438 -1381 -407 -1108
rect -334 -1181 -277 -1116
rect -334 -1208 284 -1181
rect -333 -1232 284 -1208
rect -439 -1407 -330 -1381
rect 257 -1383 281 -1232
rect 343 -1301 354 -1298
rect 257 -1388 282 -1383
rect -576 -1446 -562 -1445
rect -576 -1456 -488 -1446
rect -876 -1463 -856 -1462
rect -839 -1463 -795 -1462
rect -876 -1465 -795 -1463
rect -877 -1470 -795 -1465
rect -877 -1485 -866 -1470
rect -789 -1489 -784 -1470
rect -576 -1484 -562 -1456
rect -504 -1489 -496 -1456
rect -344 -1485 -332 -1407
rect 24 -1429 34 -1425
rect 24 -1444 132 -1429
rect 24 -1487 34 -1444
rect 96 -1493 102 -1444
rect 258 -1487 282 -1388
rect 322 -1476 330 -1436
rect 320 -1490 332 -1476
rect 343 -1493 354 -1340
rect 395 -1490 403 -1435
<< metal3 >>
rect -1311 619 -1279 1453
rect -1399 34 -1287 48
rect -1397 -427 -1378 34
rect -1347 -1 -1285 8
rect -1411 -466 -1378 -427
rect -1352 -15 -1285 -1
rect -1411 -620 -1383 -466
rect -1352 -489 -1333 -15
rect -1301 -50 -1239 -42
rect -1302 -65 -1239 -50
rect -1352 -511 -1315 -489
rect -1411 -633 -1382 -620
rect -1405 -643 -1382 -633
rect -1343 -871 -1315 -511
rect -1302 -526 -1283 -65
rect -1302 -560 -1259 -526
rect -1343 -882 -1313 -871
rect -1339 -930 -1313 -882
rect -1343 -942 -1313 -930
rect -1343 -944 -1315 -942
rect -1287 -1033 -1259 -560
rect -1290 -1115 -1259 -1033
rect -1290 -1217 -1261 -1115
rect -1297 -1255 -1252 -1217
rect -1290 -1292 -1261 -1255
rect 2 -1345 455 -1298
use PadFC  16_0
timestamp 1000338511
transform 1 0 -2500 0 1 1500
box 327 -3 1003 673
use PadFC  16_1
timestamp 1000338511
transform 0 1 1500 -1 0 2500
box 327 -3 1003 673
use PadFC  16_2
timestamp 1000338511
transform 0 -1 -1500 1 0 -2500
box 327 -3 1003 673
use PadFC  16_3
timestamp 1000338511
transform -1 0 2500 0 -1 -1500
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 1500
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 1200
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 900
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 600
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 300
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 0
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -600
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -900
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1200
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 1500 1 0 1200
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 1500 1 0 900
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 1500 1 0 600
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 1500 1 0 300
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 1500 1 0 0
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 1500 1 0 -600
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 1500 1 0 -900
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 1500 1 0 -1200
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1500
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1500
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 1500 1 0 -1500
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1500
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 1500
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1500
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 300
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 1500 -1 0 0
box -3 -11 303 1000
use top1  top1_0
timestamp 1714527017
transform 1 0 -1161 0 1 -952
box -165 -393 2536 2074
<< end >>
